magic
tech sky130A
magscale 1 2
timestamp 1640738188
<< locali >>
rect 25973 667947 26007 669341
rect 49433 668083 49467 669341
rect 63417 668151 63451 669477
rect 133889 668491 133923 669749
rect 166825 668831 166859 669953
rect 415317 668763 415351 670021
rect 427093 669851 427127 670021
rect 429209 668695 429243 669817
rect 443285 668559 443319 669817
rect 457453 668423 457487 669817
rect 471437 668355 471471 669817
rect 485789 668287 485823 669817
rect 500877 668627 500911 669817
rect 513757 668219 513791 669817
rect 527741 668015 527775 669817
rect 550005 47515 550039 47685
rect 358645 3519 358679 3689
rect 453773 3451 453807 3689
rect 361255 3417 361405 3451
rect 453589 3349 453865 3383
rect 453589 3315 453623 3349
rect 454601 2839 454635 3145
rect 582389 3043 582423 47549
<< viali >>
rect 415317 670021 415351 670055
rect 166825 669953 166859 669987
rect 133889 669749 133923 669783
rect 63417 669477 63451 669511
rect 25973 669341 26007 669375
rect 49433 669341 49467 669375
rect 166825 668797 166859 668831
rect 427093 670021 427127 670055
rect 427093 669817 427127 669851
rect 429209 669817 429243 669851
rect 415317 668729 415351 668763
rect 429209 668661 429243 668695
rect 443285 669817 443319 669851
rect 443285 668525 443319 668559
rect 457453 669817 457487 669851
rect 133889 668457 133923 668491
rect 457453 668389 457487 668423
rect 471437 669817 471471 669851
rect 471437 668321 471471 668355
rect 485789 669817 485823 669851
rect 500877 669817 500911 669851
rect 500877 668593 500911 668627
rect 513757 669817 513791 669851
rect 485789 668253 485823 668287
rect 513757 668185 513791 668219
rect 527741 669817 527775 669851
rect 63417 668117 63451 668151
rect 49433 668049 49467 668083
rect 527741 667981 527775 668015
rect 25973 667913 26007 667947
rect 550005 47685 550039 47719
rect 550005 47481 550039 47515
rect 582389 47549 582423 47583
rect 358645 3689 358679 3723
rect 358645 3485 358679 3519
rect 453773 3689 453807 3723
rect 361221 3417 361255 3451
rect 361405 3417 361439 3451
rect 453773 3417 453807 3451
rect 453865 3349 453899 3383
rect 453589 3281 453623 3315
rect 454601 3145 454635 3179
rect 582389 3009 582423 3043
rect 454601 2805 454635 2839
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 320174 700992 320180 701004
rect 154172 700964 320180 700992
rect 154172 700952 154178 700964
rect 320174 700952 320180 700964
rect 320232 700952 320238 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 316034 700924 316040 700936
rect 137888 700896 316040 700924
rect 137888 700884 137894 700896
rect 316034 700884 316040 700896
rect 316092 700884 316098 700936
rect 246942 700816 246948 700868
rect 247000 700856 247006 700868
rect 462314 700856 462320 700868
rect 247000 700828 462320 700856
rect 247000 700816 247006 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 251082 700748 251088 700800
rect 251140 700788 251146 700800
rect 478506 700788 478512 700800
rect 251140 700760 478512 700788
rect 251140 700748 251146 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 335354 700720 335360 700732
rect 89220 700692 335360 700720
rect 89220 700680 89226 700692
rect 335354 700680 335360 700692
rect 335412 700680 335418 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 329834 700652 329840 700664
rect 73028 700624 329840 700652
rect 73028 700612 73034 700624
rect 329834 700612 329840 700624
rect 329892 700612 329898 700664
rect 331858 700612 331864 700664
rect 331916 700652 331922 700664
rect 429838 700652 429844 700664
rect 331916 700624 429844 700652
rect 331916 700612 331922 700624
rect 429838 700612 429844 700624
rect 429896 700612 429902 700664
rect 233142 700544 233148 700596
rect 233200 700584 233206 700596
rect 527174 700584 527180 700596
rect 233200 700556 527180 700584
rect 233200 700544 233206 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 40494 700476 40500 700528
rect 40552 700516 40558 700528
rect 339494 700516 339500 700528
rect 40552 700488 339500 700516
rect 40552 700476 40558 700488
rect 339494 700476 339500 700488
rect 339552 700476 339558 700528
rect 170306 700408 170312 700460
rect 170364 700448 170370 700460
rect 180058 700448 180064 700460
rect 170364 700420 180064 700448
rect 170364 700408 170370 700420
rect 180058 700408 180064 700420
rect 180116 700408 180122 700460
rect 237282 700408 237288 700460
rect 237340 700448 237346 700460
rect 543458 700448 543464 700460
rect 237340 700420 543464 700448
rect 237340 700408 237346 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 349154 700380 349160 700392
rect 24360 700352 349160 700380
rect 24360 700340 24366 700352
rect 349154 700340 349160 700352
rect 349212 700340 349218 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 345014 700312 345020 700324
rect 8168 700284 345020 700312
rect 8168 700272 8174 700284
rect 345014 700272 345020 700284
rect 345072 700272 345078 700324
rect 443638 700272 443644 700324
rect 443696 700312 443702 700324
rect 494790 700312 494796 700324
rect 443696 700284 494796 700312
rect 443696 700272 443702 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 266262 700204 266268 700256
rect 266320 700244 266326 700256
rect 413646 700244 413652 700256
rect 266320 700216 413652 700244
rect 266320 700204 266326 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 260742 700136 260748 700188
rect 260800 700176 260806 700188
rect 397454 700176 397460 700188
rect 260800 700148 397460 700176
rect 260800 700136 260806 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 302234 700108 302240 700120
rect 202840 700080 302240 700108
rect 202840 700068 202846 700080
rect 302234 700068 302240 700080
rect 302292 700068 302298 700120
rect 218974 700000 218980 700052
rect 219032 700040 219038 700052
rect 306374 700040 306380 700052
rect 219032 700012 306380 700040
rect 219032 700000 219038 700012
rect 306374 700000 306380 700012
rect 306432 700000 306438 700052
rect 280062 699932 280068 699984
rect 280120 699972 280126 699984
rect 348786 699972 348792 699984
rect 280120 699944 348792 699972
rect 280120 699932 280126 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 274542 699864 274548 699916
rect 274600 699904 274606 699916
rect 332502 699904 332508 699916
rect 274600 699876 332508 699904
rect 274600 699864 274606 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 235166 699796 235172 699848
rect 235224 699836 235230 699848
rect 238018 699836 238024 699848
rect 235224 699808 238024 699836
rect 235224 699796 235230 699808
rect 238018 699796 238024 699808
rect 238076 699796 238082 699848
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 288434 699836 288440 699848
rect 267700 699808 288440 699836
rect 267700 699796 267706 699808
rect 288434 699796 288440 699808
rect 288492 699796 288498 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 292574 699768 292580 699780
rect 283892 699740 292580 699768
rect 283892 699728 283898 699740
rect 292574 699728 292580 699740
rect 292632 699728 292638 699780
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 363598 699660 363604 699712
rect 363656 699700 363662 699712
rect 364978 699700 364984 699712
rect 363656 699672 364984 699700
rect 363656 699660 363662 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 555418 699660 555424 699712
rect 555476 699700 555482 699712
rect 559650 699700 559656 699712
rect 555476 699672 559656 699700
rect 555476 699660 555482 699672
rect 559650 699660 559656 699672
rect 559708 699660 559714 699712
rect 219342 696940 219348 696992
rect 219400 696980 219406 696992
rect 580166 696980 580172 696992
rect 219400 696952 580172 696980
rect 219400 696940 219406 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 353938 683244 353944 683256
rect 3476 683216 353944 683244
rect 3476 683204 3482 683216
rect 353938 683204 353944 683216
rect 353996 683204 354002 683256
rect 223482 683136 223488 683188
rect 223540 683176 223546 683188
rect 580166 683176 580172 683188
rect 223540 683148 580172 683176
rect 223540 683136 223546 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 256602 676812 256608 676864
rect 256660 676852 256666 676864
rect 331858 676852 331864 676864
rect 256660 676824 331864 676852
rect 256660 676812 256666 676824
rect 331858 676812 331864 676824
rect 331916 676812 331922 676864
rect 283926 674500 283932 674552
rect 283984 674540 283990 674552
rect 299474 674540 299480 674552
rect 283984 674512 299480 674540
rect 283984 674500 283990 674512
rect 299474 674500 299480 674512
rect 299532 674500 299538 674552
rect 238018 674432 238024 674484
rect 238076 674472 238082 674484
rect 298002 674472 298008 674484
rect 238076 674444 298008 674472
rect 238076 674432 238082 674444
rect 298002 674432 298008 674444
rect 298060 674432 298066 674484
rect 269850 674364 269856 674416
rect 269908 674404 269914 674416
rect 363598 674404 363604 674416
rect 269908 674376 363604 674404
rect 269908 674364 269914 674376
rect 363598 674364 363604 674376
rect 363656 674364 363662 674416
rect 180058 674296 180064 674348
rect 180116 674336 180122 674348
rect 312078 674336 312084 674348
rect 180116 674308 312084 674336
rect 180116 674296 180122 674308
rect 312078 674296 312084 674308
rect 312136 674296 312142 674348
rect 241698 674228 241704 674280
rect 241756 674268 241762 674280
rect 443638 674268 443644 674280
rect 241756 674240 443644 674268
rect 241756 674228 241762 674240
rect 443638 674228 443644 674240
rect 443696 674228 443702 674280
rect 106182 674160 106188 674212
rect 106240 674200 106246 674212
rect 326154 674200 326160 674212
rect 106240 674172 326160 674200
rect 106240 674160 106246 674172
rect 326154 674160 326160 674172
rect 326212 674160 326218 674212
rect 227530 674092 227536 674144
rect 227588 674132 227594 674144
rect 555418 674132 555424 674144
rect 227588 674104 555424 674132
rect 227588 674092 227594 674104
rect 555418 674092 555424 674104
rect 555476 674092 555482 674144
rect 218146 673412 218152 673464
rect 218204 673452 218210 673464
rect 219342 673452 219348 673464
rect 218204 673424 219348 673452
rect 218204 673412 218210 673424
rect 219342 673412 219348 673424
rect 219400 673412 219406 673464
rect 232314 673412 232320 673464
rect 232372 673452 232378 673464
rect 233142 673452 233148 673464
rect 232372 673424 233148 673452
rect 232372 673412 232378 673424
rect 233142 673412 233148 673424
rect 233200 673412 233206 673464
rect 255774 673412 255780 673464
rect 255832 673452 255838 673464
rect 256602 673452 256608 673464
rect 255832 673424 256608 673452
rect 255832 673412 255838 673424
rect 256602 673412 256608 673424
rect 256660 673412 256666 673464
rect 265158 673412 265164 673464
rect 265216 673452 265222 673464
rect 266262 673452 266268 673464
rect 265216 673424 266268 673452
rect 265216 673412 265222 673424
rect 266262 673412 266268 673424
rect 266320 673412 266326 673464
rect 279234 673412 279240 673464
rect 279292 673452 279298 673464
rect 280062 673452 280068 673464
rect 279292 673424 280068 673452
rect 279292 673412 279298 673424
rect 280062 673412 280068 673424
rect 280120 673412 280126 673464
rect 204346 673344 204352 673396
rect 204404 673384 204410 673396
rect 391934 673384 391940 673396
rect 204404 673356 391940 673384
rect 204404 673344 204410 673356
rect 391934 673344 391940 673356
rect 391992 673344 391998 673396
rect 67910 673276 67916 673328
rect 67968 673316 67974 673328
rect 359458 673316 359464 673328
rect 67968 673288 359464 673316
rect 67968 673276 67974 673288
rect 359458 673276 359464 673288
rect 359516 673276 359522 673328
rect 180610 673208 180616 673260
rect 180668 673248 180674 673260
rect 555510 673248 555516 673260
rect 180668 673220 555516 673248
rect 180668 673208 180674 673220
rect 555510 673208 555516 673220
rect 555568 673208 555574 673260
rect 5166 673140 5172 673192
rect 5224 673180 5230 673192
rect 406010 673180 406016 673192
rect 5224 673152 406016 673180
rect 5224 673140 5230 673152
rect 406010 673140 406016 673152
rect 406068 673140 406074 673192
rect 5074 673072 5080 673124
rect 5132 673112 5138 673124
rect 420086 673112 420092 673124
rect 5132 673084 420092 673112
rect 5132 673072 5138 673084
rect 420086 673072 420092 673084
rect 420144 673072 420150 673124
rect 147766 673004 147772 673056
rect 147824 673044 147830 673056
rect 566642 673044 566648 673056
rect 147824 673016 566648 673044
rect 147824 673004 147830 673016
rect 566642 673004 566648 673016
rect 566700 673004 566706 673056
rect 138382 672936 138388 672988
rect 138440 672976 138446 672988
rect 576302 672976 576308 672988
rect 138440 672948 576308 672976
rect 138440 672936 138446 672948
rect 576302 672936 576308 672948
rect 576360 672936 576366 672988
rect 4982 672868 4988 672920
rect 5040 672908 5046 672920
rect 448330 672908 448336 672920
rect 5040 672880 448336 672908
rect 5040 672868 5046 672880
rect 448330 672868 448336 672880
rect 448388 672868 448394 672920
rect 124306 672800 124312 672852
rect 124364 672840 124370 672852
rect 571978 672840 571984 672852
rect 124364 672812 571984 672840
rect 124364 672800 124370 672812
rect 571978 672800 571984 672812
rect 572036 672800 572042 672852
rect 119522 672732 119528 672784
rect 119580 672772 119586 672784
rect 572070 672772 572076 672784
rect 119580 672744 572076 672772
rect 119580 672732 119586 672744
rect 572070 672732 572076 672744
rect 572128 672732 572134 672784
rect 7834 672664 7840 672716
rect 7892 672704 7898 672716
rect 462406 672704 462412 672716
rect 7892 672676 462412 672704
rect 7892 672664 7898 672676
rect 462406 672664 462412 672676
rect 462464 672664 462470 672716
rect 11882 672596 11888 672648
rect 11940 672636 11946 672648
rect 476482 672636 476488 672648
rect 11940 672608 476488 672636
rect 11940 672596 11946 672608
rect 476482 672596 476488 672608
rect 476540 672596 476546 672648
rect 105446 672528 105452 672580
rect 105504 672568 105510 672580
rect 570598 672568 570604 672580
rect 105504 672540 570604 672568
rect 105504 672528 105510 672540
rect 570598 672528 570604 672540
rect 570656 672528 570662 672580
rect 13262 672460 13268 672512
rect 13320 672500 13326 672512
rect 490558 672500 490564 672512
rect 13320 672472 490564 672500
rect 13320 672460 13326 672472
rect 490558 672460 490564 672472
rect 490616 672460 490622 672512
rect 81986 672392 81992 672444
rect 82044 672432 82050 672444
rect 558270 672432 558276 672444
rect 82044 672404 558276 672432
rect 82044 672392 82050 672404
rect 558270 672392 558276 672404
rect 558328 672392 558334 672444
rect 91370 672324 91376 672376
rect 91428 672364 91434 672376
rect 573450 672364 573456 672376
rect 91428 672336 573456 672364
rect 91428 672324 91434 672336
rect 573450 672324 573456 672336
rect 573508 672324 573514 672376
rect 96062 672256 96068 672308
rect 96120 672296 96126 672308
rect 578878 672296 578884 672308
rect 96120 672268 578884 672296
rect 96120 672256 96126 672268
rect 578878 672256 578884 672268
rect 578936 672256 578942 672308
rect 77294 672188 77300 672240
rect 77352 672228 77358 672240
rect 569310 672228 569316 672240
rect 77352 672200 569316 672228
rect 77352 672188 77358 672200
rect 569310 672188 569316 672200
rect 569368 672188 569374 672240
rect 4798 672120 4804 672172
rect 4856 672160 4862 672172
rect 499942 672160 499948 672172
rect 4856 672132 499948 672160
rect 4856 672120 4862 672132
rect 499942 672120 499948 672132
rect 500000 672120 500006 672172
rect 500862 672120 500868 672172
rect 500920 672160 500926 672172
rect 542170 672160 542176 672172
rect 500920 672132 542176 672160
rect 500920 672120 500926 672132
rect 542170 672120 542176 672132
rect 542228 672120 542234 672172
rect 7742 672052 7748 672104
rect 7800 672092 7806 672104
rect 504634 672092 504640 672104
rect 7800 672064 504640 672092
rect 7800 672052 7806 672064
rect 504634 672052 504640 672064
rect 504692 672052 504698 672104
rect 3050 671984 3056 672036
rect 3108 672024 3114 672036
rect 363782 672024 363788 672036
rect 3108 671996 363788 672024
rect 3108 671984 3114 671996
rect 363782 671984 363788 671996
rect 363840 671984 363846 672036
rect 10686 671916 10692 671968
rect 10744 671956 10750 671968
rect 373166 671956 373172 671968
rect 10744 671928 373172 671956
rect 10744 671916 10750 671928
rect 373166 671916 373172 671928
rect 373224 671916 373230 671968
rect 199378 671848 199384 671900
rect 199436 671888 199442 671900
rect 565262 671888 565268 671900
rect 199436 671860 565268 671888
rect 199436 671848 199442 671860
rect 565262 671848 565268 671860
rect 565320 671848 565326 671900
rect 213454 671780 213460 671832
rect 213512 671820 213518 671832
rect 580166 671820 580172 671832
rect 213512 671792 580172 671820
rect 213512 671780 213518 671792
rect 580166 671780 580172 671792
rect 580224 671780 580230 671832
rect 189994 671712 190000 671764
rect 190052 671752 190058 671764
rect 556982 671752 556988 671764
rect 190052 671724 556988 671752
rect 190052 671712 190058 671724
rect 556982 671712 556988 671724
rect 557040 671712 557046 671764
rect 13446 671644 13452 671696
rect 13504 671684 13510 671696
rect 401318 671684 401324 671696
rect 13504 671656 401324 671684
rect 13504 671644 13510 671656
rect 401318 671644 401324 671656
rect 401376 671644 401382 671696
rect 161842 671576 161848 671628
rect 161900 671616 161906 671628
rect 554038 671616 554044 671628
rect 161900 671588 554044 671616
rect 161900 671576 161906 671588
rect 554038 671576 554044 671588
rect 554096 671576 554102 671628
rect 12066 671508 12072 671560
rect 12124 671548 12130 671560
rect 410702 671548 410708 671560
rect 12124 671520 410708 671548
rect 12124 671508 12130 671520
rect 410702 671508 410708 671520
rect 410760 671508 410766 671560
rect 13354 671440 13360 671492
rect 13412 671480 13418 671492
rect 424778 671480 424784 671492
rect 13412 671452 424784 671480
rect 13412 671440 13418 671452
rect 424778 671440 424784 671452
rect 424836 671440 424842 671492
rect 143074 671372 143080 671424
rect 143132 671412 143138 671424
rect 561030 671412 561036 671424
rect 143132 671384 561036 671412
rect 143132 671372 143138 671384
rect 561030 671372 561036 671384
rect 561088 671372 561094 671424
rect 7926 671304 7932 671356
rect 7984 671344 7990 671356
rect 438854 671344 438860 671356
rect 7984 671316 438860 671344
rect 7984 671304 7990 671316
rect 438854 671304 438860 671316
rect 438912 671304 438918 671356
rect 9030 671236 9036 671288
rect 9088 671276 9094 671288
rect 453022 671276 453028 671288
rect 9088 671248 453028 671276
rect 9088 671236 9094 671248
rect 453022 671236 453028 671248
rect 453080 671236 453086 671288
rect 114830 671168 114836 671220
rect 114888 671208 114894 671220
rect 565170 671208 565176 671220
rect 114888 671180 565176 671208
rect 114888 671168 114894 671180
rect 565170 671168 565176 671180
rect 565228 671168 565234 671220
rect 10410 671100 10416 671152
rect 10468 671140 10474 671152
rect 467098 671140 467104 671152
rect 10468 671112 467104 671140
rect 10468 671100 10474 671112
rect 467098 671100 467104 671112
rect 467156 671100 467162 671152
rect 11790 671032 11796 671084
rect 11848 671072 11854 671084
rect 481174 671072 481180 671084
rect 11848 671044 481180 671072
rect 11848 671032 11854 671044
rect 481174 671032 481180 671044
rect 481232 671032 481238 671084
rect 86678 670964 86684 671016
rect 86736 671004 86742 671016
rect 555418 671004 555424 671016
rect 86736 670976 555424 671004
rect 86736 670964 86742 670976
rect 555418 670964 555424 670976
rect 555476 670964 555482 671016
rect 13170 670896 13176 670948
rect 13228 670936 13234 670948
rect 495250 670936 495256 670948
rect 13228 670908 495256 670936
rect 13228 670896 13234 670908
rect 495250 670896 495256 670908
rect 495308 670896 495314 670948
rect 7650 670828 7656 670880
rect 7708 670868 7714 670880
rect 509326 670868 509332 670880
rect 7708 670840 509332 670868
rect 7708 670828 7714 670840
rect 509326 670828 509332 670840
rect 509384 670828 509390 670880
rect 58526 670760 58532 670812
rect 58584 670800 58590 670812
rect 573358 670800 573364 670812
rect 58584 670772 573364 670800
rect 58584 670760 58590 670772
rect 573358 670760 573364 670772
rect 573416 670760 573422 670812
rect 44450 670692 44456 670744
rect 44508 670732 44514 670744
rect 569218 670732 569224 670744
rect 44508 670704 569224 670732
rect 44508 670692 44514 670704
rect 569218 670692 569224 670704
rect 569276 670692 569282 670744
rect 6362 670624 6368 670676
rect 6420 670664 6426 670676
rect 359090 670664 359096 670676
rect 6420 670636 359096 670664
rect 6420 670624 6426 670636
rect 359090 670624 359096 670636
rect 359148 670624 359154 670676
rect 359458 670624 359464 670676
rect 359516 670664 359522 670676
rect 580350 670664 580356 670676
rect 359516 670636 580356 670664
rect 359516 670624 359522 670636
rect 580350 670624 580356 670636
rect 580408 670624 580414 670676
rect 8018 670556 8024 670608
rect 8076 670596 8082 670608
rect 368474 670596 368480 670608
rect 8076 670568 368480 670596
rect 8076 670556 8082 670568
rect 368474 670556 368480 670568
rect 368532 670556 368538 670608
rect 204070 670488 204076 670540
rect 204128 670528 204134 670540
rect 566734 670528 566740 670540
rect 204128 670500 566740 670528
rect 204128 670488 204134 670500
rect 566734 670488 566740 670500
rect 566792 670488 566798 670540
rect 3878 670420 3884 670472
rect 3936 670460 3942 670472
rect 204346 670460 204352 670472
rect 3936 670432 204352 670460
rect 3936 670420 3942 670432
rect 204346 670420 204352 670432
rect 204404 670420 204410 670472
rect 208762 670420 208768 670472
rect 208820 670460 208826 670472
rect 574922 670460 574928 670472
rect 208820 670432 574928 670460
rect 208820 670420 208826 670432
rect 574922 670420 574928 670432
rect 574980 670420 574986 670472
rect 9214 670352 9220 670404
rect 9272 670392 9278 670404
rect 377858 670392 377864 670404
rect 9272 670364 377864 670392
rect 9272 670352 9278 670364
rect 377858 670352 377864 670364
rect 377916 670352 377922 670404
rect 9122 670284 9128 670336
rect 9180 670324 9186 670336
rect 382550 670324 382556 670336
rect 9180 670296 382556 670324
rect 9180 670284 9186 670296
rect 382550 670284 382556 670296
rect 382608 670284 382614 670336
rect 12158 670216 12164 670268
rect 12216 670256 12222 670268
rect 387242 670256 387248 670268
rect 12216 670228 387248 670256
rect 12216 670216 12222 670228
rect 387242 670216 387248 670228
rect 387300 670216 387306 670268
rect 185302 670148 185308 670200
rect 185360 670188 185366 670200
rect 562502 670188 562508 670200
rect 185360 670160 562508 670188
rect 185360 670148 185366 670160
rect 562502 670148 562508 670160
rect 562560 670148 562566 670200
rect 175918 670080 175924 670132
rect 175976 670120 175982 670132
rect 555602 670120 555608 670132
rect 175976 670092 555608 670120
rect 175976 670080 175982 670092
rect 555602 670080 555608 670092
rect 555660 670080 555666 670132
rect 10594 670012 10600 670064
rect 10652 670052 10658 670064
rect 396350 670052 396356 670064
rect 10652 670024 396356 670052
rect 10652 670012 10658 670024
rect 396350 670012 396356 670024
rect 396408 670012 396414 670064
rect 415302 670052 415308 670064
rect 415263 670024 415308 670052
rect 415302 670012 415308 670024
rect 415360 670012 415366 670064
rect 427081 670055 427139 670061
rect 427081 670021 427093 670055
rect 427127 670052 427139 670055
rect 433886 670052 433892 670064
rect 427127 670024 433892 670052
rect 427127 670021 427139 670024
rect 427081 670015 427139 670021
rect 433886 670012 433892 670024
rect 433944 670012 433950 670064
rect 166810 669984 166816 669996
rect 166771 669956 166816 669984
rect 166810 669944 166816 669956
rect 166868 669944 166874 669996
rect 171594 669944 171600 669996
rect 171652 669984 171658 669996
rect 561122 669984 561128 669996
rect 171652 669956 561128 669984
rect 171652 669944 171658 669956
rect 561122 669944 561128 669956
rect 561180 669944 561186 669996
rect 157058 669876 157064 669928
rect 157116 669916 157122 669928
rect 558362 669916 558368 669928
rect 157116 669888 558368 669916
rect 157116 669876 157122 669888
rect 558362 669876 558368 669888
rect 558420 669876 558426 669928
rect 11974 669808 11980 669860
rect 12032 669848 12038 669860
rect 427081 669851 427139 669857
rect 427081 669848 427093 669851
rect 12032 669820 427093 669848
rect 12032 669808 12038 669820
rect 427081 669817 427093 669820
rect 427127 669817 427139 669851
rect 429194 669848 429200 669860
rect 429155 669820 429200 669848
rect 427081 669811 427139 669817
rect 429194 669808 429200 669820
rect 429252 669808 429258 669860
rect 443270 669848 443276 669860
rect 443231 669820 443276 669848
rect 443270 669808 443276 669820
rect 443328 669808 443334 669860
rect 457438 669848 457444 669860
rect 457399 669820 457444 669848
rect 457438 669808 457444 669820
rect 457496 669808 457502 669860
rect 471422 669848 471428 669860
rect 471383 669820 471428 669848
rect 471422 669808 471428 669820
rect 471480 669808 471486 669860
rect 485774 669848 485780 669860
rect 485735 669820 485780 669848
rect 485774 669808 485780 669820
rect 485832 669808 485838 669860
rect 500862 669848 500868 669860
rect 500823 669820 500868 669848
rect 500862 669808 500868 669820
rect 500920 669808 500926 669860
rect 513742 669848 513748 669860
rect 513703 669820 513748 669848
rect 513742 669808 513748 669820
rect 513800 669808 513806 669860
rect 527726 669848 527732 669860
rect 527687 669820 527732 669848
rect 527726 669808 527732 669820
rect 527784 669808 527790 669860
rect 133874 669780 133880 669792
rect 133835 669752 133880 669780
rect 133874 669740 133880 669752
rect 133932 669740 133938 669792
rect 152826 669740 152832 669792
rect 152884 669780 152890 669792
rect 580442 669780 580448 669792
rect 152884 669752 580448 669780
rect 152884 669740 152890 669752
rect 580442 669740 580448 669752
rect 580500 669740 580506 669792
rect 129274 669672 129280 669724
rect 129332 669712 129338 669724
rect 562410 669712 562416 669724
rect 129332 669684 562416 669712
rect 129332 669672 129338 669684
rect 562410 669672 562416 669684
rect 562468 669672 562474 669724
rect 110322 669604 110328 669656
rect 110380 669644 110386 669656
rect 566550 669644 566556 669656
rect 110380 669616 566556 669644
rect 110380 669604 110386 669616
rect 566550 669604 566556 669616
rect 566608 669604 566614 669656
rect 101122 669536 101128 669588
rect 101180 669576 101186 669588
rect 576210 669576 576216 669588
rect 101180 669548 576216 669576
rect 101180 669536 101186 669548
rect 576210 669536 576216 669548
rect 576268 669536 576274 669588
rect 63402 669508 63408 669520
rect 63363 669480 63408 669508
rect 63402 669468 63408 669480
rect 63460 669468 63466 669520
rect 72970 669468 72976 669520
rect 73028 669508 73034 669520
rect 574830 669508 574836 669520
rect 73028 669480 574836 669508
rect 73028 669468 73034 669480
rect 574830 669468 574836 669480
rect 574888 669468 574894 669520
rect 39942 669400 39948 669452
rect 40000 669440 40006 669452
rect 560938 669440 560944 669452
rect 40000 669412 560944 669440
rect 40000 669400 40006 669412
rect 560938 669400 560944 669412
rect 560996 669400 561002 669452
rect 25958 669372 25964 669384
rect 25919 669344 25964 669372
rect 25958 669332 25964 669344
rect 26016 669332 26022 669384
rect 49418 669372 49424 669384
rect 49379 669344 49424 669372
rect 49418 669332 49424 669344
rect 49476 669332 49482 669384
rect 54202 669332 54208 669384
rect 54260 669372 54266 669384
rect 580258 669372 580264 669384
rect 54260 669344 580264 669372
rect 54260 669332 54266 669344
rect 580258 669332 580264 669344
rect 580316 669332 580322 669384
rect 194686 669196 194692 669248
rect 194744 669236 194750 669248
rect 194744 669208 200114 669236
rect 194744 669196 194750 669208
rect 200086 668896 200114 669208
rect 554130 668896 554136 668908
rect 200086 668868 554136 668896
rect 554130 668856 554136 668868
rect 554188 668856 554194 668908
rect 166813 668831 166871 668837
rect 166813 668797 166825 668831
rect 166859 668828 166871 668831
rect 556890 668828 556896 668840
rect 166859 668800 556896 668828
rect 166859 668797 166871 668800
rect 166813 668791 166871 668797
rect 556890 668788 556896 668800
rect 556948 668788 556954 668840
rect 6270 668720 6276 668772
rect 6328 668760 6334 668772
rect 415305 668763 415363 668769
rect 415305 668760 415317 668763
rect 6328 668732 415317 668760
rect 6328 668720 6334 668732
rect 415305 668729 415317 668732
rect 415351 668729 415363 668763
rect 415305 668723 415363 668729
rect 3786 668652 3792 668704
rect 3844 668692 3850 668704
rect 429197 668695 429255 668701
rect 429197 668692 429209 668695
rect 3844 668664 429209 668692
rect 3844 668652 3850 668664
rect 429197 668661 429209 668664
rect 429243 668661 429255 668695
rect 429197 668655 429255 668661
rect 3418 668584 3424 668636
rect 3476 668624 3482 668636
rect 500865 668627 500923 668633
rect 500865 668624 500877 668627
rect 3476 668596 500877 668624
rect 3476 668584 3482 668596
rect 500865 668593 500877 668596
rect 500911 668593 500923 668627
rect 500865 668587 500923 668593
rect 10502 668516 10508 668568
rect 10560 668556 10566 668568
rect 443273 668559 443331 668565
rect 443273 668556 443285 668559
rect 10560 668528 443285 668556
rect 10560 668516 10566 668528
rect 443273 668525 443285 668528
rect 443319 668525 443331 668559
rect 443273 668519 443331 668525
rect 133877 668491 133935 668497
rect 133877 668457 133889 668491
rect 133923 668488 133935 668491
rect 578970 668488 578976 668500
rect 133923 668460 578976 668488
rect 133923 668457 133935 668460
rect 133877 668451 133935 668457
rect 578970 668448 578976 668460
rect 579028 668448 579034 668500
rect 3694 668380 3700 668432
rect 3752 668420 3758 668432
rect 457441 668423 457499 668429
rect 457441 668420 457453 668423
rect 3752 668392 457453 668420
rect 3752 668380 3758 668392
rect 457441 668389 457453 668392
rect 457487 668389 457499 668423
rect 457441 668383 457499 668389
rect 4890 668312 4896 668364
rect 4948 668352 4954 668364
rect 471425 668355 471483 668361
rect 471425 668352 471437 668355
rect 4948 668324 471437 668352
rect 4948 668312 4954 668324
rect 471425 668321 471437 668324
rect 471471 668321 471483 668355
rect 471425 668315 471483 668321
rect 3602 668244 3608 668296
rect 3660 668284 3666 668296
rect 485777 668287 485835 668293
rect 485777 668284 485789 668287
rect 3660 668256 485789 668284
rect 3660 668244 3666 668256
rect 485777 668253 485789 668256
rect 485823 668253 485835 668287
rect 485777 668247 485835 668253
rect 3510 668176 3516 668228
rect 3568 668216 3574 668228
rect 513745 668219 513803 668225
rect 513745 668216 513757 668219
rect 3568 668188 513757 668216
rect 3568 668176 3574 668188
rect 513745 668185 513757 668188
rect 513791 668185 513803 668219
rect 513745 668179 513803 668185
rect 63405 668151 63463 668157
rect 63405 668117 63417 668151
rect 63451 668148 63463 668151
rect 574738 668148 574744 668160
rect 63451 668120 574744 668148
rect 63451 668117 63463 668120
rect 63405 668111 63463 668117
rect 574738 668108 574744 668120
rect 574796 668108 574802 668160
rect 49421 668083 49479 668089
rect 49421 668049 49433 668083
rect 49467 668080 49479 668083
rect 565078 668080 565084 668092
rect 49467 668052 565084 668080
rect 49467 668049 49479 668052
rect 49421 668043 49479 668049
rect 565078 668040 565084 668052
rect 565136 668040 565142 668092
rect 7558 667972 7564 668024
rect 7616 668012 7622 668024
rect 527729 668015 527787 668021
rect 527729 668012 527741 668015
rect 7616 667984 527741 668012
rect 7616 667972 7622 667984
rect 527729 667981 527741 667984
rect 527775 667981 527787 668015
rect 527729 667975 527787 667981
rect 25961 667947 26019 667953
rect 25961 667913 25973 667947
rect 26007 667944 26019 667947
rect 562318 667944 562324 667956
rect 26007 667916 562324 667944
rect 26007 667913 26019 667916
rect 25961 667907 26019 667913
rect 562318 667904 562324 667916
rect 562376 667904 562382 667956
rect 3234 658180 3240 658232
rect 3292 658220 3298 658232
rect 6362 658220 6368 658232
rect 3292 658192 6368 658220
rect 3292 658180 3298 658192
rect 6362 658180 6368 658192
rect 6420 658180 6426 658232
rect 566734 644376 566740 644428
rect 566792 644416 566798 644428
rect 580166 644416 580172 644428
rect 566792 644388 580172 644416
rect 566792 644376 566798 644388
rect 580166 644376 580172 644388
rect 580224 644376 580230 644428
rect 3326 632136 3332 632188
rect 3384 632176 3390 632188
rect 8018 632176 8024 632188
rect 3384 632148 8024 632176
rect 3384 632136 3390 632148
rect 8018 632136 8024 632148
rect 8076 632136 8082 632188
rect 574922 632000 574928 632052
rect 574980 632040 574986 632052
rect 579706 632040 579712 632052
rect 574980 632012 579712 632040
rect 574980 632000 574986 632012
rect 579706 632000 579712 632012
rect 579764 632000 579770 632052
rect 2958 619284 2964 619336
rect 3016 619324 3022 619336
rect 9214 619324 9220 619336
rect 3016 619296 9220 619324
rect 3016 619284 3022 619296
rect 9214 619284 9220 619296
rect 9272 619284 9278 619336
rect 565262 618196 565268 618248
rect 565320 618236 565326 618248
rect 579798 618236 579804 618248
rect 565320 618208 579804 618236
rect 565320 618196 565326 618208
rect 579798 618196 579804 618208
rect 579856 618196 579862 618248
rect 2866 607112 2872 607164
rect 2924 607152 2930 607164
rect 10686 607152 10692 607164
rect 2924 607124 10692 607152
rect 2924 607112 2930 607124
rect 10686 607112 10692 607124
rect 10744 607112 10750 607164
rect 556982 591948 556988 592000
rect 557040 591988 557046 592000
rect 580166 591988 580172 592000
rect 557040 591960 580172 591988
rect 557040 591948 557046 591960
rect 580166 591948 580172 591960
rect 580224 591948 580230 592000
rect 3142 580456 3148 580508
rect 3200 580496 3206 580508
rect 9122 580496 9128 580508
rect 3200 580468 9128 580496
rect 3200 580456 3206 580468
rect 9122 580456 9128 580468
rect 9180 580456 9186 580508
rect 554130 578144 554136 578196
rect 554188 578184 554194 578196
rect 580166 578184 580172 578196
rect 554188 578156 580172 578184
rect 554188 578144 554194 578156
rect 580166 578144 580172 578156
rect 580224 578144 580230 578196
rect 562502 564340 562508 564392
rect 562560 564380 562566 564392
rect 580166 564380 580172 564392
rect 562560 564352 580172 564380
rect 562560 564340 562566 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 3326 554684 3332 554736
rect 3384 554724 3390 554736
rect 12158 554724 12164 554736
rect 3384 554696 12164 554724
rect 3384 554684 3390 554696
rect 12158 554684 12164 554696
rect 12216 554684 12222 554736
rect 555602 538160 555608 538212
rect 555660 538200 555666 538212
rect 580166 538200 580172 538212
rect 555660 538172 580172 538200
rect 555660 538160 555666 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 3234 528504 3240 528556
rect 3292 528544 3298 528556
rect 10594 528544 10600 528556
rect 3292 528516 10600 528544
rect 3292 528504 3298 528516
rect 10594 528504 10600 528516
rect 10652 528504 10658 528556
rect 555510 525716 555516 525768
rect 555568 525756 555574 525768
rect 580166 525756 580172 525768
rect 555568 525728 580172 525756
rect 555568 525716 555574 525728
rect 580166 525716 580172 525728
rect 580224 525716 580230 525768
rect 2774 515584 2780 515636
rect 2832 515624 2838 515636
rect 5166 515624 5172 515636
rect 2832 515596 5172 515624
rect 2832 515584 2838 515596
rect 5166 515584 5172 515596
rect 5224 515584 5230 515636
rect 561122 511912 561128 511964
rect 561180 511952 561186 511964
rect 580166 511952 580172 511964
rect 561180 511924 580172 511952
rect 561180 511912 561186 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 3326 502256 3332 502308
rect 3384 502296 3390 502308
rect 13446 502296 13452 502308
rect 3384 502268 13452 502296
rect 3384 502256 3390 502268
rect 13446 502256 13452 502268
rect 13504 502256 13510 502308
rect 554038 485732 554044 485784
rect 554096 485772 554102 485784
rect 580166 485772 580172 485784
rect 554096 485744 580172 485772
rect 554096 485732 554102 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 3326 476008 3332 476060
rect 3384 476048 3390 476060
rect 12066 476048 12072 476060
rect 3384 476020 12072 476048
rect 3384 476008 3390 476020
rect 12066 476008 12072 476020
rect 12124 476008 12130 476060
rect 556890 471928 556896 471980
rect 556948 471968 556954 471980
rect 580166 471968 580172 471980
rect 556948 471940 580172 471968
rect 556948 471928 556954 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 2774 463428 2780 463480
rect 2832 463468 2838 463480
rect 5074 463468 5080 463480
rect 2832 463440 5080 463468
rect 2832 463428 2838 463440
rect 5074 463428 5080 463440
rect 5132 463428 5138 463480
rect 558362 458124 558368 458176
rect 558420 458164 558426 458176
rect 580166 458164 580172 458176
rect 558420 458136 580172 458164
rect 558420 458124 558426 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 2958 449556 2964 449608
rect 3016 449596 3022 449608
rect 6270 449596 6276 449608
rect 3016 449568 6276 449596
rect 3016 449556 3022 449568
rect 6270 449556 6276 449568
rect 6328 449556 6334 449608
rect 566642 431876 566648 431928
rect 566700 431916 566706 431928
rect 580166 431916 580172 431928
rect 566700 431888 580172 431916
rect 566700 431876 566706 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 13354 423620 13360 423632
rect 3384 423592 13360 423620
rect 3384 423580 3390 423592
rect 13354 423580 13360 423592
rect 13412 423580 13418 423632
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 11974 411244 11980 411256
rect 3384 411216 11980 411244
rect 3384 411204 3390 411216
rect 11974 411204 11980 411216
rect 12032 411204 12038 411256
rect 561030 405628 561036 405680
rect 561088 405668 561094 405680
rect 580166 405668 580172 405680
rect 561088 405640 580172 405668
rect 561088 405628 561094 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 3326 371560 3332 371612
rect 3384 371600 3390 371612
rect 7926 371600 7932 371612
rect 3384 371572 7932 371600
rect 3384 371560 3390 371572
rect 7926 371560 7932 371572
rect 7984 371560 7990 371612
rect 576302 365644 576308 365696
rect 576360 365684 576366 365696
rect 579982 365684 579988 365696
rect 576360 365656 579988 365684
rect 576360 365644 576366 365656
rect 579982 365644 579988 365656
rect 580040 365644 580046 365696
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 4982 358476 4988 358488
rect 2832 358448 4988 358476
rect 2832 358436 2838 358448
rect 4982 358436 4988 358448
rect 5040 358436 5046 358488
rect 562410 353200 562416 353252
rect 562468 353240 562474 353252
rect 580166 353240 580172 353252
rect 562468 353212 580172 353240
rect 562468 353200 562474 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 2958 346332 2964 346384
rect 3016 346372 3022 346384
rect 10502 346372 10508 346384
rect 3016 346344 10508 346372
rect 3016 346332 3022 346344
rect 10502 346332 10508 346344
rect 10560 346332 10566 346384
rect 572070 325592 572076 325644
rect 572128 325632 572134 325644
rect 580166 325632 580172 325644
rect 572128 325604 580172 325632
rect 572128 325592 572134 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3234 320016 3240 320068
rect 3292 320056 3298 320068
rect 9030 320056 9036 320068
rect 3292 320028 9036 320056
rect 3292 320016 3298 320028
rect 9030 320016 9036 320028
rect 9088 320016 9094 320068
rect 571978 313216 571984 313268
rect 572036 313256 572042 313268
rect 580166 313256 580172 313268
rect 572036 313228 580172 313256
rect 572036 313216 572042 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3326 306212 3332 306264
rect 3384 306252 3390 306264
rect 7834 306252 7840 306264
rect 3384 306224 7840 306252
rect 3384 306212 3390 306224
rect 7834 306212 7840 306224
rect 7892 306212 7898 306264
rect 565170 299412 565176 299464
rect 565228 299452 565234 299464
rect 580166 299452 580172 299464
rect 565228 299424 580172 299452
rect 565228 299412 565234 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 570598 273164 570604 273216
rect 570656 273204 570662 273216
rect 580166 273204 580172 273216
rect 570656 273176 580172 273204
rect 570656 273164 570662 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3234 267656 3240 267708
rect 3292 267696 3298 267708
rect 10410 267696 10416 267708
rect 3292 267668 10416 267696
rect 3292 267656 3298 267668
rect 10410 267656 10416 267668
rect 10468 267656 10474 267708
rect 566550 259360 566556 259412
rect 566608 259400 566614 259412
rect 579614 259400 579620 259412
rect 566608 259372 579620 259400
rect 566608 259360 566614 259372
rect 579614 259360 579620 259372
rect 579672 259360 579678 259412
rect 3326 255212 3332 255264
rect 3384 255252 3390 255264
rect 11882 255252 11888 255264
rect 3384 255224 11888 255252
rect 3384 255212 3390 255224
rect 11882 255212 11888 255224
rect 11940 255212 11946 255264
rect 576210 245556 576216 245608
rect 576268 245596 576274 245608
rect 580166 245596 580172 245608
rect 576268 245568 580172 245596
rect 576268 245556 576274 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 2774 241068 2780 241120
rect 2832 241108 2838 241120
rect 4890 241108 4896 241120
rect 2832 241080 4896 241108
rect 2832 241068 2838 241080
rect 4890 241068 4896 241080
rect 4948 241068 4954 241120
rect 573450 233180 573456 233232
rect 573508 233220 573514 233232
rect 580166 233220 580172 233232
rect 573508 233192 580172 233220
rect 573508 233180 573514 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 11790 215268 11796 215280
rect 3384 215240 11796 215268
rect 3384 215228 3390 215240
rect 11790 215228 11796 215240
rect 11848 215228 11854 215280
rect 555418 206932 555424 206984
rect 555476 206972 555482 206984
rect 579890 206972 579896 206984
rect 555476 206944 579896 206972
rect 555476 206932 555482 206944
rect 579890 206932 579896 206944
rect 579948 206932 579954 206984
rect 3326 202784 3332 202836
rect 3384 202824 3390 202836
rect 13262 202824 13268 202836
rect 3384 202796 13268 202824
rect 3384 202784 3390 202796
rect 13262 202784 13268 202796
rect 13320 202784 13326 202836
rect 569310 193128 569316 193180
rect 569368 193168 569374 193180
rect 580166 193168 580172 193180
rect 569368 193140 580172 193168
rect 569368 193128 569374 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 558270 179324 558276 179376
rect 558328 179364 558334 179376
rect 580166 179364 580172 179376
rect 558328 179336 580172 179364
rect 558328 179324 558334 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 574830 166948 574836 167000
rect 574888 166988 574894 167000
rect 580166 166988 580172 167000
rect 574888 166960 580172 166988
rect 574888 166948 574894 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 13170 164200 13176 164212
rect 3384 164172 13176 164200
rect 3384 164160 3390 164172
rect 13170 164160 13176 164172
rect 13228 164160 13234 164212
rect 574738 153144 574744 153196
rect 574796 153184 574802 153196
rect 579614 153184 579620 153196
rect 574796 153156 579620 153184
rect 574796 153144 574802 153156
rect 579614 153144 579620 153156
rect 579672 153144 579678 153196
rect 3602 150356 3608 150408
rect 3660 150396 3666 150408
rect 7742 150396 7748 150408
rect 3660 150368 7748 150396
rect 3660 150356 3666 150368
rect 7742 150356 7748 150368
rect 7800 150356 7806 150408
rect 2774 136824 2780 136876
rect 2832 136864 2838 136876
rect 4798 136864 4804 136876
rect 2832 136836 4804 136864
rect 2832 136824 2838 136836
rect 4798 136824 4804 136836
rect 4856 136824 4862 136876
rect 573358 126896 573364 126948
rect 573416 126936 573422 126948
rect 580166 126936 580172 126948
rect 573416 126908 580172 126936
rect 573416 126896 573422 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 565078 113092 565084 113144
rect 565136 113132 565142 113144
rect 580166 113132 580172 113144
rect 565136 113104 580172 113132
rect 565136 113092 565142 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 2958 111120 2964 111172
rect 3016 111160 3022 111172
rect 7650 111160 7656 111172
rect 3016 111132 7656 111160
rect 3016 111120 3022 111132
rect 7650 111120 7656 111132
rect 7708 111120 7714 111172
rect 3234 97928 3240 97980
rect 3292 97968 3298 97980
rect 11698 97968 11704 97980
rect 3292 97940 11704 97968
rect 3292 97928 3298 97940
rect 11698 97928 11704 97940
rect 11756 97928 11762 97980
rect 569218 86912 569224 86964
rect 569276 86952 569282 86964
rect 580166 86952 580172 86964
rect 569276 86924 580172 86952
rect 569276 86912 569282 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 576118 73108 576124 73160
rect 576176 73148 576182 73160
rect 580166 73148 580172 73160
rect 576176 73120 580172 73148
rect 576176 73108 576182 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3510 71612 3516 71664
rect 3568 71652 3574 71664
rect 8938 71652 8944 71664
rect 3568 71624 8944 71652
rect 3568 71612 3574 71624
rect 8938 71612 8944 71624
rect 8996 71612 9002 71664
rect 560938 60664 560944 60716
rect 560996 60704 561002 60716
rect 580166 60704 580172 60716
rect 560996 60676 580172 60704
rect 560996 60664 561002 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 13078 59344 13084 59356
rect 3108 59316 13084 59344
rect 3108 59304 3114 59316
rect 13078 59304 13084 59316
rect 13136 59304 13142 59356
rect 171134 48288 171140 48340
rect 171192 48288 171198 48340
rect 12250 48220 12256 48272
rect 12308 48260 12314 48272
rect 24302 48260 24308 48272
rect 12308 48232 24308 48260
rect 12308 48220 12314 48232
rect 24302 48220 24308 48232
rect 24360 48220 24366 48272
rect 27430 48220 27436 48272
rect 27488 48260 27494 48272
rect 38470 48260 38476 48272
rect 27488 48232 38476 48260
rect 27488 48220 27494 48232
rect 38470 48220 38476 48232
rect 38528 48220 38534 48272
rect 45462 48220 45468 48272
rect 45520 48260 45526 48272
rect 54938 48260 54944 48272
rect 45520 48232 54944 48260
rect 45520 48220 45526 48232
rect 54938 48220 54944 48232
rect 54996 48220 55002 48272
rect 171152 48260 171180 48288
rect 172146 48260 172152 48272
rect 171152 48232 172152 48260
rect 172146 48220 172152 48232
rect 172204 48220 172210 48272
rect 4062 48152 4068 48204
rect 4120 48192 4126 48204
rect 16574 48192 16580 48204
rect 4120 48164 16580 48192
rect 4120 48152 4126 48164
rect 16574 48152 16580 48164
rect 16632 48152 16638 48204
rect 17862 48152 17868 48204
rect 17920 48192 17926 48204
rect 29730 48192 29736 48204
rect 17920 48164 29736 48192
rect 17920 48152 17926 48164
rect 29730 48152 29736 48164
rect 29788 48152 29794 48204
rect 33042 48152 33048 48204
rect 33100 48192 33106 48204
rect 43990 48192 43996 48204
rect 33100 48164 43996 48192
rect 33100 48152 33106 48164
rect 43990 48152 43996 48164
rect 44048 48152 44054 48204
rect 48222 48152 48228 48204
rect 48280 48192 48286 48204
rect 58250 48192 58256 48204
rect 48280 48164 58256 48192
rect 48280 48152 48286 48164
rect 58250 48152 58256 48164
rect 58308 48152 58314 48204
rect 59262 48152 59268 48204
rect 59320 48192 59326 48204
rect 68094 48192 68100 48204
rect 59320 48164 68100 48192
rect 59320 48152 59326 48164
rect 68094 48152 68100 48164
rect 68152 48152 68158 48204
rect 73062 48152 73068 48204
rect 73120 48192 73126 48204
rect 81250 48192 81256 48204
rect 73120 48164 81256 48192
rect 73120 48152 73126 48164
rect 81250 48152 81256 48164
rect 81308 48152 81314 48204
rect 8202 48084 8208 48136
rect 8260 48124 8266 48136
rect 20990 48124 20996 48136
rect 8260 48096 20996 48124
rect 8260 48084 8266 48096
rect 20990 48084 20996 48096
rect 21048 48084 21054 48136
rect 24762 48084 24768 48136
rect 24820 48124 24826 48136
rect 36354 48124 36360 48136
rect 24820 48096 36360 48124
rect 24820 48084 24826 48096
rect 36354 48084 36360 48096
rect 36412 48084 36418 48136
rect 41322 48084 41328 48136
rect 41380 48124 41386 48136
rect 51626 48124 51632 48136
rect 41380 48096 51632 48124
rect 41380 48084 41386 48096
rect 51626 48084 51632 48096
rect 51684 48084 51690 48136
rect 52362 48084 52368 48136
rect 52420 48124 52426 48136
rect 61470 48124 61476 48136
rect 52420 48096 61476 48124
rect 52420 48084 52426 48096
rect 61470 48084 61476 48096
rect 61528 48084 61534 48136
rect 67542 48084 67548 48136
rect 67600 48124 67606 48136
rect 75730 48124 75736 48136
rect 67600 48096 75736 48124
rect 67600 48084 67606 48096
rect 75730 48084 75736 48096
rect 75788 48084 75794 48136
rect 95050 48084 95056 48136
rect 95108 48124 95114 48136
rect 102042 48124 102048 48136
rect 95108 48096 102048 48124
rect 95108 48084 95114 48096
rect 102042 48084 102048 48096
rect 102100 48084 102106 48136
rect 12342 48016 12348 48068
rect 12400 48056 12406 48068
rect 25406 48056 25412 48068
rect 12400 48028 25412 48056
rect 12400 48016 12406 48028
rect 25406 48016 25412 48028
rect 25464 48016 25470 48068
rect 28902 48016 28908 48068
rect 28960 48056 28966 48068
rect 39574 48056 39580 48068
rect 28960 48028 39580 48056
rect 28960 48016 28966 48028
rect 39574 48016 39580 48028
rect 39632 48016 39638 48068
rect 39942 48016 39948 48068
rect 40000 48056 40006 48068
rect 50522 48056 50528 48068
rect 40000 48028 50528 48056
rect 40000 48016 40006 48028
rect 50522 48016 50528 48028
rect 50580 48016 50586 48068
rect 50982 48016 50988 48068
rect 51040 48056 51046 48068
rect 60458 48056 60464 48068
rect 51040 48028 60464 48056
rect 51040 48016 51046 48028
rect 60458 48016 60464 48028
rect 60516 48016 60522 48068
rect 61930 48016 61936 48068
rect 61988 48056 61994 48068
rect 70302 48056 70308 48068
rect 61988 48028 70308 48056
rect 61988 48016 61994 48028
rect 70302 48016 70308 48028
rect 70360 48016 70366 48068
rect 77938 48056 77944 48068
rect 71516 48028 77944 48056
rect 13722 47948 13728 48000
rect 13780 47988 13786 48000
rect 26418 47988 26424 48000
rect 13780 47960 26424 47988
rect 13780 47948 13786 47960
rect 26418 47948 26424 47960
rect 26476 47948 26482 48000
rect 30282 47948 30288 48000
rect 30340 47988 30346 48000
rect 41782 47988 41788 48000
rect 30340 47960 41788 47988
rect 30340 47948 30346 47960
rect 41782 47948 41788 47960
rect 41840 47948 41846 48000
rect 42702 47948 42708 48000
rect 42760 47988 42766 48000
rect 52730 47988 52736 48000
rect 42760 47960 52736 47988
rect 42760 47948 42766 47960
rect 52730 47948 52736 47960
rect 52788 47948 52794 48000
rect 62022 47948 62028 48000
rect 62080 47988 62086 48000
rect 71406 47988 71412 48000
rect 62080 47960 71412 47988
rect 62080 47948 62086 47960
rect 71406 47948 71412 47960
rect 71464 47948 71470 48000
rect 6822 47880 6828 47932
rect 6880 47920 6886 47932
rect 19886 47920 19892 47932
rect 6880 47892 19892 47920
rect 6880 47880 6886 47892
rect 19886 47880 19892 47892
rect 19944 47880 19950 47932
rect 26142 47880 26148 47932
rect 26200 47920 26206 47932
rect 37458 47920 37464 47932
rect 26200 47892 37464 47920
rect 26200 47880 26206 47892
rect 37458 47880 37464 47892
rect 37516 47880 37522 47932
rect 38562 47880 38568 47932
rect 38620 47920 38626 47932
rect 49510 47920 49516 47932
rect 38620 47892 49516 47920
rect 38620 47880 38626 47892
rect 49510 47880 49516 47892
rect 49568 47880 49574 47932
rect 53650 47880 53656 47932
rect 53708 47920 53714 47932
rect 62574 47920 62580 47932
rect 53708 47892 62580 47920
rect 53708 47880 53714 47892
rect 62574 47880 62580 47892
rect 62632 47880 62638 47932
rect 63402 47880 63408 47932
rect 63460 47920 63466 47932
rect 63460 47892 68692 47920
rect 63460 47880 63466 47892
rect 5442 47812 5448 47864
rect 5500 47852 5506 47864
rect 18782 47852 18788 47864
rect 5500 47824 18788 47852
rect 5500 47812 5506 47824
rect 18782 47812 18788 47824
rect 18840 47812 18846 47864
rect 19242 47812 19248 47864
rect 19300 47852 19306 47864
rect 30834 47852 30840 47864
rect 19300 47824 30840 47852
rect 19300 47812 19306 47824
rect 30834 47812 30840 47824
rect 30892 47812 30898 47864
rect 31662 47812 31668 47864
rect 31720 47852 31726 47864
rect 42886 47852 42892 47864
rect 31720 47824 42892 47852
rect 31720 47812 31726 47824
rect 42886 47812 42892 47824
rect 42944 47812 42950 47864
rect 44082 47812 44088 47864
rect 44140 47852 44146 47864
rect 53834 47852 53840 47864
rect 44140 47824 53840 47852
rect 44140 47812 44146 47824
rect 53834 47812 53840 47824
rect 53892 47812 53898 47864
rect 55122 47812 55128 47864
rect 55180 47852 55186 47864
rect 64782 47852 64788 47864
rect 55180 47824 64788 47852
rect 55180 47812 55186 47824
rect 64782 47812 64788 47824
rect 64840 47812 64846 47864
rect 68664 47852 68692 47892
rect 70302 47880 70308 47932
rect 70360 47920 70366 47932
rect 71516 47920 71544 48028
rect 77938 48016 77944 48028
rect 77996 48016 78002 48068
rect 79962 48016 79968 48068
rect 80020 48056 80026 48068
rect 87782 48056 87788 48068
rect 80020 48028 87788 48056
rect 80020 48016 80026 48028
rect 87782 48016 87788 48028
rect 87840 48016 87846 48068
rect 91002 48016 91008 48068
rect 91060 48056 91066 48068
rect 97626 48056 97632 48068
rect 91060 48028 97632 48056
rect 91060 48016 91066 48028
rect 97626 48016 97632 48028
rect 97684 48016 97690 48068
rect 92382 47948 92388 48000
rect 92440 47988 92446 48000
rect 98730 47988 98736 48000
rect 92440 47960 98736 47988
rect 92440 47948 92446 47960
rect 98730 47948 98736 47960
rect 98788 47948 98794 48000
rect 102042 47948 102048 48000
rect 102100 47988 102106 48000
rect 107562 47988 107568 48000
rect 102100 47960 107568 47988
rect 102100 47948 102106 47960
rect 107562 47948 107568 47960
rect 107620 47948 107626 48000
rect 531406 47948 531412 48000
rect 531464 47988 531470 48000
rect 531464 47960 536880 47988
rect 531464 47948 531470 47960
rect 70360 47892 71544 47920
rect 70360 47880 70366 47892
rect 74442 47880 74448 47932
rect 74500 47920 74506 47932
rect 82354 47920 82360 47932
rect 74500 47892 82360 47920
rect 74500 47880 74506 47892
rect 82354 47880 82360 47892
rect 82412 47880 82418 47932
rect 86770 47880 86776 47932
rect 86828 47920 86834 47932
rect 93302 47920 93308 47932
rect 86828 47892 93308 47920
rect 86828 47880 86834 47892
rect 93302 47880 93308 47892
rect 93360 47880 93366 47932
rect 103330 47880 103336 47932
rect 103388 47920 103394 47932
rect 108574 47920 108580 47932
rect 103388 47892 108580 47920
rect 103388 47880 103394 47892
rect 108574 47880 108580 47892
rect 108632 47880 108638 47932
rect 115842 47880 115848 47932
rect 115900 47920 115906 47932
rect 120626 47920 120632 47932
rect 115900 47892 120632 47920
rect 115900 47880 115906 47892
rect 120626 47880 120632 47892
rect 120684 47880 120690 47932
rect 135162 47880 135168 47932
rect 135220 47920 135226 47932
rect 138198 47920 138204 47932
rect 135220 47892 138204 47920
rect 135220 47880 135226 47892
rect 138198 47880 138204 47892
rect 138256 47880 138262 47932
rect 146202 47880 146208 47932
rect 146260 47920 146266 47932
rect 149146 47920 149152 47932
rect 146260 47892 149152 47920
rect 146260 47880 146266 47892
rect 149146 47880 149152 47892
rect 149204 47880 149210 47932
rect 158622 47880 158628 47932
rect 158680 47920 158686 47932
rect 160094 47920 160100 47932
rect 158680 47892 160100 47920
rect 158680 47880 158686 47892
rect 160094 47880 160100 47892
rect 160152 47880 160158 47932
rect 212718 47880 212724 47932
rect 212776 47920 212782 47932
rect 214006 47920 214012 47932
rect 212776 47892 214012 47920
rect 212776 47880 212782 47892
rect 214006 47880 214012 47892
rect 214064 47880 214070 47932
rect 536852 47920 536880 47960
rect 536926 47948 536932 48000
rect 536984 47988 536990 48000
rect 538122 47988 538128 48000
rect 536984 47960 538128 47988
rect 536984 47948 536990 47960
rect 538122 47948 538128 47960
rect 538180 47948 538186 48000
rect 546770 47948 546776 48000
rect 546828 47988 546834 48000
rect 547782 47988 547788 48000
rect 546828 47960 547788 47988
rect 546828 47948 546834 47960
rect 547782 47948 547788 47960
rect 547840 47948 547846 48000
rect 547874 47948 547880 48000
rect 547932 47988 547938 48000
rect 549070 47988 549076 48000
rect 547932 47960 549076 47988
rect 547932 47948 547938 47960
rect 549070 47948 549076 47960
rect 549128 47948 549134 48000
rect 557534 47920 557540 47932
rect 536852 47892 557540 47920
rect 557534 47880 557540 47892
rect 557592 47880 557598 47932
rect 72510 47852 72516 47864
rect 68664 47824 72516 47852
rect 72510 47812 72516 47824
rect 72568 47812 72574 47864
rect 74626 47852 74632 47864
rect 74506 47824 74632 47852
rect 2682 47744 2688 47796
rect 2740 47784 2746 47796
rect 15470 47784 15476 47796
rect 2740 47756 15476 47784
rect 2740 47744 2746 47756
rect 15470 47744 15476 47756
rect 15528 47744 15534 47796
rect 20622 47744 20628 47796
rect 20680 47784 20686 47796
rect 31938 47784 31944 47796
rect 20680 47756 31944 47784
rect 20680 47744 20686 47756
rect 31938 47744 31944 47756
rect 31996 47744 32002 47796
rect 35802 47744 35808 47796
rect 35860 47784 35866 47796
rect 46198 47784 46204 47796
rect 35860 47756 46204 47784
rect 35860 47744 35866 47756
rect 46198 47744 46204 47756
rect 46256 47744 46262 47796
rect 46842 47744 46848 47796
rect 46900 47784 46906 47796
rect 57146 47784 57152 47796
rect 46900 47756 57152 47784
rect 46900 47744 46906 47756
rect 57146 47744 57152 47756
rect 57204 47744 57210 47796
rect 57882 47744 57888 47796
rect 57940 47784 57946 47796
rect 66990 47784 66996 47796
rect 57940 47756 66996 47784
rect 57940 47744 57946 47756
rect 66990 47744 66996 47756
rect 67048 47744 67054 47796
rect 9582 47676 9588 47728
rect 9640 47716 9646 47728
rect 22094 47716 22100 47728
rect 9640 47688 22100 47716
rect 9640 47676 9646 47688
rect 22094 47676 22100 47688
rect 22152 47676 22158 47728
rect 23382 47676 23388 47728
rect 23440 47716 23446 47728
rect 35250 47716 35256 47728
rect 23440 47688 35256 47716
rect 23440 47676 23446 47688
rect 35250 47676 35256 47688
rect 35308 47676 35314 47728
rect 37090 47676 37096 47728
rect 37148 47716 37154 47728
rect 47302 47716 47308 47728
rect 37148 47688 47308 47716
rect 37148 47676 37154 47688
rect 47302 47676 47308 47688
rect 47360 47676 47366 47728
rect 53742 47676 53748 47728
rect 53800 47716 53806 47728
rect 63678 47716 63684 47728
rect 53800 47688 63684 47716
rect 53800 47676 53806 47688
rect 63678 47676 63684 47688
rect 63736 47676 63742 47728
rect 64782 47676 64788 47728
rect 64840 47716 64846 47728
rect 64840 47688 66116 47716
rect 64840 47676 64846 47688
rect 3970 47608 3976 47660
rect 4028 47648 4034 47660
rect 17678 47648 17684 47660
rect 4028 47620 17684 47648
rect 4028 47608 4034 47620
rect 17678 47608 17684 47620
rect 17736 47608 17742 47660
rect 28810 47608 28816 47660
rect 28868 47648 28874 47660
rect 40678 47648 40684 47660
rect 28868 47620 40684 47648
rect 28868 47608 28874 47620
rect 40678 47608 40684 47620
rect 40736 47608 40742 47660
rect 45370 47608 45376 47660
rect 45428 47648 45434 47660
rect 56042 47648 56048 47660
rect 45428 47620 56048 47648
rect 45428 47608 45434 47620
rect 56042 47608 56048 47620
rect 56100 47608 56106 47660
rect 56502 47608 56508 47660
rect 56560 47648 56566 47660
rect 65886 47648 65892 47660
rect 56560 47620 65892 47648
rect 56560 47608 56566 47620
rect 65886 47608 65892 47620
rect 65944 47608 65950 47660
rect 66088 47648 66116 47688
rect 66162 47676 66168 47728
rect 66220 47716 66226 47728
rect 74506 47716 74534 47824
rect 74626 47812 74632 47824
rect 74684 47812 74690 47864
rect 84102 47812 84108 47864
rect 84160 47852 84166 47864
rect 91094 47852 91100 47864
rect 84160 47824 91100 47852
rect 84160 47812 84166 47824
rect 91094 47812 91100 47824
rect 91152 47812 91158 47864
rect 93762 47812 93768 47864
rect 93820 47852 93826 47864
rect 99834 47852 99840 47864
rect 93820 47824 99840 47852
rect 93820 47812 93826 47824
rect 99834 47812 99840 47824
rect 99892 47812 99898 47864
rect 107562 47812 107568 47864
rect 107620 47852 107626 47864
rect 112990 47852 112996 47864
rect 107620 47824 112996 47852
rect 107620 47812 107626 47824
rect 112990 47812 112996 47824
rect 113048 47812 113054 47864
rect 114462 47812 114468 47864
rect 114520 47852 114526 47864
rect 119614 47852 119620 47864
rect 114520 47824 119620 47852
rect 114520 47812 114526 47824
rect 119614 47812 119620 47824
rect 119672 47812 119678 47864
rect 130378 47812 130384 47864
rect 130436 47852 130442 47864
rect 131666 47852 131672 47864
rect 130436 47824 131672 47852
rect 130436 47812 130442 47824
rect 131666 47812 131672 47824
rect 131724 47812 131730 47864
rect 137278 47812 137284 47864
rect 137336 47852 137342 47864
rect 140406 47852 140412 47864
rect 137336 47824 140412 47852
rect 137336 47812 137342 47824
rect 140406 47812 140412 47824
rect 140464 47812 140470 47864
rect 144822 47812 144828 47864
rect 144880 47852 144886 47864
rect 146938 47852 146944 47864
rect 144880 47824 146944 47852
rect 144880 47812 144886 47824
rect 146938 47812 146944 47824
rect 146996 47812 147002 47864
rect 148962 47812 148968 47864
rect 149020 47852 149026 47864
rect 151354 47852 151360 47864
rect 149020 47824 151360 47852
rect 149020 47812 149026 47824
rect 151354 47812 151360 47824
rect 151412 47812 151418 47864
rect 153102 47812 153108 47864
rect 153160 47852 153166 47864
rect 154666 47852 154672 47864
rect 153160 47824 154672 47852
rect 153160 47812 153166 47824
rect 154666 47812 154672 47824
rect 154724 47812 154730 47864
rect 155862 47812 155868 47864
rect 155920 47852 155926 47864
rect 157886 47852 157892 47864
rect 155920 47824 157892 47852
rect 155920 47812 155926 47824
rect 157886 47812 157892 47824
rect 157944 47812 157950 47864
rect 160002 47812 160008 47864
rect 160060 47852 160066 47864
rect 161198 47852 161204 47864
rect 160060 47824 161204 47852
rect 160060 47812 160066 47824
rect 161198 47812 161204 47824
rect 161256 47812 161262 47864
rect 162762 47812 162768 47864
rect 162820 47852 162826 47864
rect 164510 47852 164516 47864
rect 162820 47824 164516 47852
rect 162820 47812 162826 47824
rect 164510 47812 164516 47824
rect 164568 47812 164574 47864
rect 166902 47812 166908 47864
rect 166960 47852 166966 47864
rect 167730 47852 167736 47864
rect 166960 47824 167736 47852
rect 166960 47812 166966 47824
rect 167730 47812 167736 47824
rect 167788 47812 167794 47864
rect 176654 47812 176660 47864
rect 176712 47852 176718 47864
rect 177666 47852 177672 47864
rect 176712 47824 177672 47852
rect 176712 47812 176718 47824
rect 177666 47812 177672 47824
rect 177724 47812 177730 47864
rect 186314 47812 186320 47864
rect 186372 47852 186378 47864
rect 187510 47852 187516 47864
rect 186372 47824 187516 47852
rect 186372 47812 186378 47824
rect 187510 47812 187516 47824
rect 187568 47812 187574 47864
rect 206094 47812 206100 47864
rect 206152 47852 206158 47864
rect 206922 47852 206928 47864
rect 206152 47824 206928 47852
rect 206152 47812 206158 47824
rect 206922 47812 206928 47824
rect 206980 47812 206986 47864
rect 217042 47812 217048 47864
rect 217100 47852 217106 47864
rect 217962 47852 217968 47864
rect 217100 47824 217968 47852
rect 217100 47812 217106 47824
rect 217962 47812 217968 47824
rect 218020 47812 218026 47864
rect 222562 47812 222568 47864
rect 222620 47852 222626 47864
rect 223482 47852 223488 47864
rect 222620 47824 223488 47852
rect 222620 47812 222626 47824
rect 223482 47812 223488 47824
rect 223540 47812 223546 47864
rect 226886 47812 226892 47864
rect 226944 47852 226950 47864
rect 227622 47852 227628 47864
rect 226944 47824 227628 47852
rect 226944 47812 226950 47824
rect 227622 47812 227628 47824
rect 227680 47812 227686 47864
rect 227990 47812 227996 47864
rect 228048 47852 228054 47864
rect 229002 47852 229008 47864
rect 228048 47824 229008 47852
rect 228048 47812 228054 47824
rect 229002 47812 229008 47824
rect 229060 47812 229066 47864
rect 229094 47812 229100 47864
rect 229152 47852 229158 47864
rect 231946 47852 231952 47864
rect 229152 47824 231952 47852
rect 229152 47812 229158 47824
rect 231946 47812 231952 47824
rect 232004 47812 232010 47864
rect 232406 47812 232412 47864
rect 232464 47852 232470 47864
rect 233142 47852 233148 47864
rect 232464 47824 233148 47852
rect 232464 47812 232470 47824
rect 233142 47812 233148 47824
rect 233200 47812 233206 47864
rect 233510 47812 233516 47864
rect 233568 47852 233574 47864
rect 234522 47852 234528 47864
rect 233568 47824 234528 47852
rect 233568 47812 233574 47824
rect 234522 47812 234528 47824
rect 234580 47812 234586 47864
rect 234614 47812 234620 47864
rect 234672 47852 234678 47864
rect 237466 47852 237472 47864
rect 234672 47824 237472 47852
rect 234672 47812 234678 47824
rect 237466 47812 237472 47824
rect 237524 47812 237530 47864
rect 237834 47812 237840 47864
rect 237892 47852 237898 47864
rect 238662 47852 238668 47864
rect 237892 47824 238668 47852
rect 237892 47812 237898 47824
rect 238662 47812 238668 47824
rect 238720 47812 238726 47864
rect 240042 47812 240048 47864
rect 240100 47852 240106 47864
rect 240778 47852 240784 47864
rect 240100 47824 240784 47852
rect 240100 47812 240106 47824
rect 240778 47812 240784 47824
rect 240836 47812 240842 47864
rect 244458 47812 244464 47864
rect 244516 47852 244522 47864
rect 245562 47852 245568 47864
rect 244516 47824 245568 47852
rect 244516 47812 244522 47824
rect 245562 47812 245568 47824
rect 245620 47812 245626 47864
rect 248874 47812 248880 47864
rect 248932 47852 248938 47864
rect 249702 47852 249708 47864
rect 248932 47824 249708 47852
rect 248932 47812 248938 47824
rect 249702 47812 249708 47824
rect 249760 47812 249766 47864
rect 249886 47812 249892 47864
rect 249944 47852 249950 47864
rect 250990 47852 250996 47864
rect 249944 47824 250996 47852
rect 249944 47812 249950 47824
rect 250990 47812 250996 47824
rect 251048 47812 251054 47864
rect 254302 47812 254308 47864
rect 254360 47852 254366 47864
rect 255222 47852 255228 47864
rect 254360 47824 255228 47852
rect 254360 47812 254366 47824
rect 255222 47812 255228 47824
rect 255280 47812 255286 47864
rect 255406 47812 255412 47864
rect 255464 47852 255470 47864
rect 256510 47852 256516 47864
rect 255464 47824 256516 47852
rect 255464 47812 255470 47824
rect 256510 47812 256516 47824
rect 256568 47812 256574 47864
rect 260926 47812 260932 47864
rect 260984 47852 260990 47864
rect 264238 47852 264244 47864
rect 260984 47824 264244 47852
rect 260984 47812 260990 47824
rect 264238 47812 264244 47824
rect 264296 47812 264302 47864
rect 270770 47812 270776 47864
rect 270828 47852 270834 47864
rect 271782 47852 271788 47864
rect 270828 47824 271788 47852
rect 270828 47812 270834 47824
rect 271782 47812 271788 47824
rect 271840 47812 271846 47864
rect 281718 47812 281724 47864
rect 281776 47852 281782 47864
rect 282730 47852 282736 47864
rect 281776 47824 282736 47852
rect 281776 47812 281782 47824
rect 282730 47812 282736 47824
rect 282788 47812 282794 47864
rect 286042 47812 286048 47864
rect 286100 47852 286106 47864
rect 286962 47852 286968 47864
rect 286100 47824 286968 47852
rect 286100 47812 286106 47824
rect 286962 47812 286968 47824
rect 287020 47812 287026 47864
rect 287146 47812 287152 47864
rect 287204 47852 287210 47864
rect 288342 47852 288348 47864
rect 287204 47824 288348 47852
rect 287204 47812 287210 47824
rect 288342 47812 288348 47824
rect 288400 47812 288406 47864
rect 291562 47812 291568 47864
rect 291620 47852 291626 47864
rect 292482 47852 292488 47864
rect 291620 47824 292488 47852
rect 291620 47812 291626 47824
rect 292482 47812 292488 47824
rect 292540 47812 292546 47864
rect 292666 47812 292672 47864
rect 292724 47852 292730 47864
rect 293770 47852 293776 47864
rect 292724 47824 293776 47852
rect 292724 47812 292730 47824
rect 293770 47812 293776 47824
rect 293828 47812 293834 47864
rect 296990 47812 296996 47864
rect 297048 47852 297054 47864
rect 298002 47852 298008 47864
rect 297048 47824 298008 47852
rect 297048 47812 297054 47824
rect 298002 47812 298008 47824
rect 298060 47812 298066 47864
rect 301406 47812 301412 47864
rect 301464 47852 301470 47864
rect 302142 47852 302148 47864
rect 301464 47824 302148 47852
rect 301464 47812 301470 47824
rect 302142 47812 302148 47824
rect 302200 47812 302206 47864
rect 302510 47812 302516 47864
rect 302568 47852 302574 47864
rect 303522 47852 303528 47864
rect 302568 47824 303528 47852
rect 302568 47812 302574 47824
rect 303522 47812 303528 47824
rect 303580 47812 303586 47864
rect 303614 47812 303620 47864
rect 303672 47852 303678 47864
rect 304902 47852 304908 47864
rect 303672 47824 304908 47852
rect 303672 47812 303678 47824
rect 304902 47812 304908 47824
rect 304960 47812 304966 47864
rect 307938 47812 307944 47864
rect 307996 47852 308002 47864
rect 308950 47852 308956 47864
rect 307996 47824 308956 47852
rect 307996 47812 308002 47824
rect 308950 47812 308956 47824
rect 309008 47812 309014 47864
rect 312354 47812 312360 47864
rect 312412 47852 312418 47864
rect 313182 47852 313188 47864
rect 312412 47824 313188 47852
rect 312412 47812 312418 47824
rect 313182 47812 313188 47824
rect 313240 47812 313246 47864
rect 317874 47812 317880 47864
rect 317932 47852 317938 47864
rect 318702 47852 318708 47864
rect 317932 47824 318708 47852
rect 317932 47812 317938 47824
rect 318702 47812 318708 47824
rect 318760 47812 318766 47864
rect 324406 47812 324412 47864
rect 324464 47852 324470 47864
rect 325510 47852 325516 47864
rect 324464 47824 325516 47852
rect 324464 47812 324470 47824
rect 325510 47812 325516 47824
rect 325568 47812 325574 47864
rect 328822 47812 328828 47864
rect 328880 47852 328886 47864
rect 329742 47852 329748 47864
rect 328880 47824 329748 47852
rect 328880 47812 328886 47824
rect 329742 47812 329748 47824
rect 329800 47812 329806 47864
rect 329926 47812 329932 47864
rect 329984 47852 329990 47864
rect 331122 47852 331128 47864
rect 329984 47824 331128 47852
rect 329984 47812 329990 47824
rect 331122 47812 331128 47824
rect 331180 47812 331186 47864
rect 334250 47812 334256 47864
rect 334308 47852 334314 47864
rect 335262 47852 335268 47864
rect 334308 47824 335268 47852
rect 334308 47812 334314 47824
rect 335262 47812 335268 47824
rect 335320 47812 335326 47864
rect 335354 47812 335360 47864
rect 335412 47852 335418 47864
rect 336642 47852 336648 47864
rect 335412 47824 336648 47852
rect 335412 47812 335418 47824
rect 336642 47812 336648 47824
rect 336700 47812 336706 47864
rect 339770 47812 339776 47864
rect 339828 47852 339834 47864
rect 340782 47852 340788 47864
rect 339828 47824 340788 47852
rect 339828 47812 339834 47824
rect 340782 47812 340788 47824
rect 340840 47812 340846 47864
rect 350718 47812 350724 47864
rect 350776 47852 350782 47864
rect 351730 47852 351736 47864
rect 350776 47824 351736 47852
rect 350776 47812 350782 47824
rect 351730 47812 351736 47824
rect 351788 47812 351794 47864
rect 355042 47812 355048 47864
rect 355100 47852 355106 47864
rect 355962 47852 355968 47864
rect 355100 47824 355968 47852
rect 355100 47812 355106 47824
rect 355962 47812 355968 47824
rect 356020 47812 356026 47864
rect 360562 47812 360568 47864
rect 360620 47852 360626 47864
rect 361482 47852 361488 47864
rect 360620 47824 361488 47852
rect 360620 47812 360626 47824
rect 361482 47812 361488 47824
rect 361540 47812 361546 47864
rect 366082 47812 366088 47864
rect 366140 47852 366146 47864
rect 367002 47852 367008 47864
rect 366140 47824 367008 47852
rect 366140 47812 366146 47824
rect 367002 47812 367008 47824
rect 367060 47812 367066 47864
rect 367094 47812 367100 47864
rect 367152 47852 367158 47864
rect 368290 47852 368296 47864
rect 367152 47824 368296 47852
rect 367152 47812 367158 47824
rect 368290 47812 368296 47824
rect 368348 47812 368354 47864
rect 371510 47812 371516 47864
rect 371568 47852 371574 47864
rect 372522 47852 372528 47864
rect 371568 47824 372528 47852
rect 371568 47812 371574 47824
rect 372522 47812 372528 47824
rect 372580 47812 372586 47864
rect 372614 47812 372620 47864
rect 372672 47852 372678 47864
rect 373810 47852 373816 47864
rect 372672 47824 373816 47852
rect 372672 47812 372678 47824
rect 373810 47812 373816 47824
rect 373868 47812 373874 47864
rect 375926 47812 375932 47864
rect 375984 47852 375990 47864
rect 376662 47852 376668 47864
rect 375984 47824 376668 47852
rect 375984 47812 375990 47824
rect 376662 47812 376668 47824
rect 376720 47812 376726 47864
rect 377030 47812 377036 47864
rect 377088 47852 377094 47864
rect 378042 47852 378048 47864
rect 377088 47824 378048 47852
rect 377088 47812 377094 47824
rect 378042 47812 378048 47824
rect 378100 47812 378106 47864
rect 378134 47812 378140 47864
rect 378192 47852 378198 47864
rect 379422 47852 379428 47864
rect 378192 47824 379428 47852
rect 378192 47812 378198 47824
rect 379422 47812 379428 47824
rect 379480 47812 379486 47864
rect 382458 47812 382464 47864
rect 382516 47852 382522 47864
rect 383470 47852 383476 47864
rect 382516 47824 383476 47852
rect 382516 47812 382522 47824
rect 383470 47812 383476 47824
rect 383528 47812 383534 47864
rect 386874 47812 386880 47864
rect 386932 47852 386938 47864
rect 387702 47852 387708 47864
rect 386932 47824 387708 47852
rect 386932 47812 386938 47824
rect 387702 47812 387708 47824
rect 387760 47812 387766 47864
rect 387978 47812 387984 47864
rect 388036 47852 388042 47864
rect 389082 47852 389088 47864
rect 388036 47824 389088 47852
rect 388036 47812 388042 47824
rect 389082 47812 389088 47824
rect 389140 47812 389146 47864
rect 392302 47812 392308 47864
rect 392360 47852 392366 47864
rect 393222 47852 393228 47864
rect 392360 47824 393228 47852
rect 392360 47812 392366 47824
rect 393222 47812 393228 47824
rect 393280 47812 393286 47864
rect 403250 47812 403256 47864
rect 403308 47852 403314 47864
rect 404262 47852 404268 47864
rect 403308 47824 404268 47852
rect 403308 47812 403314 47824
rect 404262 47812 404268 47824
rect 404320 47812 404326 47864
rect 404354 47812 404360 47864
rect 404412 47852 404418 47864
rect 405642 47852 405648 47864
rect 404412 47824 405648 47852
rect 404412 47812 404418 47824
rect 405642 47812 405648 47824
rect 405700 47812 405706 47864
rect 408770 47812 408776 47864
rect 408828 47852 408834 47864
rect 409782 47852 409788 47864
rect 408828 47824 409788 47852
rect 408828 47812 408834 47824
rect 409782 47812 409788 47824
rect 409840 47812 409846 47864
rect 409874 47812 409880 47864
rect 409932 47852 409938 47864
rect 411070 47852 411076 47864
rect 409932 47824 411076 47852
rect 409932 47812 409938 47824
rect 411070 47812 411076 47824
rect 411128 47812 411134 47864
rect 418614 47812 418620 47864
rect 418672 47852 418678 47864
rect 419442 47852 419448 47864
rect 418672 47824 419448 47852
rect 418672 47812 418678 47824
rect 419442 47812 419448 47824
rect 419500 47812 419506 47864
rect 419718 47812 419724 47864
rect 419776 47852 419782 47864
rect 420730 47852 420736 47864
rect 419776 47824 420736 47852
rect 419776 47812 419782 47824
rect 420730 47812 420736 47824
rect 420788 47812 420794 47864
rect 429562 47812 429568 47864
rect 429620 47852 429626 47864
rect 430482 47852 430488 47864
rect 429620 47824 430488 47852
rect 429620 47812 429626 47824
rect 430482 47812 430488 47824
rect 430540 47812 430546 47864
rect 430666 47812 430672 47864
rect 430724 47852 430730 47864
rect 431862 47852 431868 47864
rect 430724 47824 431868 47852
rect 430724 47812 430730 47824
rect 431862 47812 431868 47824
rect 431920 47812 431926 47864
rect 436186 47812 436192 47864
rect 436244 47852 436250 47864
rect 437290 47852 437296 47864
rect 436244 47824 437296 47852
rect 436244 47812 436250 47824
rect 437290 47812 437296 47824
rect 437348 47812 437354 47864
rect 439406 47812 439412 47864
rect 439464 47852 439470 47864
rect 440142 47852 440148 47864
rect 439464 47824 440148 47852
rect 439464 47812 439470 47824
rect 440142 47812 440148 47824
rect 440200 47812 440206 47864
rect 440510 47812 440516 47864
rect 440568 47852 440574 47864
rect 441522 47852 441528 47864
rect 440568 47824 441528 47852
rect 440568 47812 440574 47824
rect 441522 47812 441528 47824
rect 441580 47812 441586 47864
rect 441614 47812 441620 47864
rect 441672 47852 441678 47864
rect 442902 47852 442908 47864
rect 441672 47824 442908 47852
rect 441672 47812 441678 47824
rect 442902 47812 442908 47824
rect 442960 47812 442966 47864
rect 446030 47812 446036 47864
rect 446088 47852 446094 47864
rect 447042 47852 447048 47864
rect 446088 47824 447048 47852
rect 446088 47812 446094 47824
rect 447042 47812 447048 47824
rect 447100 47812 447106 47864
rect 450354 47812 450360 47864
rect 450412 47852 450418 47864
rect 451182 47852 451188 47864
rect 450412 47824 451188 47852
rect 450412 47812 450418 47824
rect 451182 47812 451188 47824
rect 451240 47812 451246 47864
rect 451458 47812 451464 47864
rect 451516 47852 451522 47864
rect 452562 47852 452568 47864
rect 451516 47824 452568 47852
rect 451516 47812 451522 47824
rect 452562 47812 452568 47824
rect 452620 47812 452626 47864
rect 456978 47812 456984 47864
rect 457036 47852 457042 47864
rect 457990 47852 457996 47864
rect 457036 47824 457996 47852
rect 457036 47812 457042 47824
rect 457990 47812 457996 47824
rect 458048 47812 458054 47864
rect 461302 47812 461308 47864
rect 461360 47852 461366 47864
rect 462222 47852 462228 47864
rect 461360 47824 462228 47852
rect 461360 47812 461366 47824
rect 462222 47812 462228 47824
rect 462280 47812 462286 47864
rect 466822 47812 466828 47864
rect 466880 47852 466886 47864
rect 467742 47852 467748 47864
rect 466880 47824 467748 47852
rect 466880 47812 466886 47824
rect 467742 47812 467748 47824
rect 467800 47812 467806 47864
rect 467926 47812 467932 47864
rect 467984 47852 467990 47864
rect 469122 47852 469128 47864
rect 467984 47824 469128 47852
rect 467984 47812 467990 47824
rect 469122 47812 469128 47824
rect 469180 47812 469186 47864
rect 472250 47812 472256 47864
rect 472308 47852 472314 47864
rect 473262 47852 473268 47864
rect 472308 47824 473268 47852
rect 472308 47812 472314 47824
rect 473262 47812 473268 47824
rect 473320 47812 473326 47864
rect 473354 47812 473360 47864
rect 473412 47852 473418 47864
rect 474550 47852 474556 47864
rect 473412 47824 474556 47852
rect 473412 47812 473418 47824
rect 474550 47812 474556 47824
rect 474608 47812 474614 47864
rect 477770 47812 477776 47864
rect 477828 47852 477834 47864
rect 478782 47852 478788 47864
rect 477828 47824 478788 47852
rect 477828 47812 477834 47824
rect 478782 47812 478788 47824
rect 478840 47812 478846 47864
rect 478874 47812 478880 47864
rect 478932 47852 478938 47864
rect 480070 47852 480076 47864
rect 478932 47824 480076 47852
rect 478932 47812 478938 47824
rect 480070 47812 480076 47824
rect 480128 47812 480134 47864
rect 483290 47812 483296 47864
rect 483348 47852 483354 47864
rect 484210 47852 484216 47864
rect 483348 47824 484216 47852
rect 483348 47812 483354 47824
rect 484210 47812 484216 47824
rect 484268 47812 484274 47864
rect 493134 47812 493140 47864
rect 493192 47852 493198 47864
rect 493962 47852 493968 47864
rect 493192 47824 493968 47852
rect 493192 47812 493198 47824
rect 493962 47812 493968 47824
rect 494020 47812 494026 47864
rect 494238 47812 494244 47864
rect 494296 47852 494302 47864
rect 495342 47852 495348 47864
rect 494296 47824 495348 47852
rect 494296 47812 494302 47824
rect 495342 47812 495348 47824
rect 495400 47812 495406 47864
rect 499666 47812 499672 47864
rect 499724 47852 499730 47864
rect 500770 47852 500776 47864
rect 499724 47824 500776 47852
rect 499724 47812 499730 47824
rect 500770 47812 500776 47824
rect 500828 47812 500834 47864
rect 504082 47812 504088 47864
rect 504140 47852 504146 47864
rect 505002 47852 505008 47864
rect 504140 47824 505008 47852
rect 504140 47812 504146 47824
rect 505002 47812 505008 47824
rect 505060 47812 505066 47864
rect 508406 47812 508412 47864
rect 508464 47852 508470 47864
rect 509142 47852 509148 47864
rect 508464 47824 509148 47852
rect 508464 47812 508470 47824
rect 509142 47812 509148 47824
rect 509200 47812 509206 47864
rect 510614 47812 510620 47864
rect 510672 47852 510678 47864
rect 511902 47852 511908 47864
rect 510672 47824 511908 47852
rect 510672 47812 510678 47824
rect 511902 47812 511908 47824
rect 511960 47812 511966 47864
rect 513926 47812 513932 47864
rect 513984 47852 513990 47864
rect 514662 47852 514668 47864
rect 513984 47824 514668 47852
rect 513984 47812 513990 47824
rect 514662 47812 514668 47824
rect 514720 47812 514726 47864
rect 515030 47812 515036 47864
rect 515088 47852 515094 47864
rect 516042 47852 516048 47864
rect 515088 47824 516048 47852
rect 515088 47812 515094 47824
rect 516042 47812 516048 47824
rect 516100 47812 516106 47864
rect 516134 47812 516140 47864
rect 516192 47852 516198 47864
rect 517422 47852 517428 47864
rect 516192 47824 517428 47852
rect 516192 47812 516198 47824
rect 517422 47812 517428 47824
rect 517480 47812 517486 47864
rect 519354 47812 519360 47864
rect 519412 47852 519418 47864
rect 520182 47852 520188 47864
rect 519412 47824 520188 47852
rect 519412 47812 519418 47824
rect 520182 47812 520188 47824
rect 520240 47812 520246 47864
rect 520458 47812 520464 47864
rect 520516 47852 520522 47864
rect 521562 47852 521568 47864
rect 520516 47824 521568 47852
rect 520516 47812 520522 47824
rect 521562 47812 521568 47824
rect 521620 47812 521626 47864
rect 524874 47812 524880 47864
rect 524932 47852 524938 47864
rect 525702 47852 525708 47864
rect 524932 47824 525708 47852
rect 524932 47812 524938 47824
rect 525702 47812 525708 47824
rect 525760 47812 525766 47864
rect 525978 47812 525984 47864
rect 526036 47852 526042 47864
rect 526990 47852 526996 47864
rect 526036 47824 526996 47852
rect 526036 47812 526042 47824
rect 526990 47812 526996 47824
rect 527048 47812 527054 47864
rect 530394 47812 530400 47864
rect 530452 47852 530458 47864
rect 531222 47852 531228 47864
rect 530452 47824 531228 47852
rect 530452 47812 530458 47824
rect 531222 47812 531228 47824
rect 531280 47812 531286 47864
rect 535822 47812 535828 47864
rect 535880 47852 535886 47864
rect 536742 47852 536748 47864
rect 535880 47824 536748 47852
rect 535880 47812 535886 47824
rect 536742 47812 536748 47824
rect 536800 47812 536806 47864
rect 560938 47852 560944 47864
rect 536944 47824 560944 47852
rect 77202 47744 77208 47796
rect 77260 47784 77266 47796
rect 84562 47784 84568 47796
rect 77260 47756 84568 47784
rect 77260 47744 77266 47756
rect 84562 47744 84568 47756
rect 84620 47744 84626 47796
rect 86862 47744 86868 47796
rect 86920 47784 86926 47796
rect 94406 47784 94412 47796
rect 86920 47756 94412 47784
rect 86920 47744 86926 47756
rect 94406 47744 94412 47756
rect 94464 47744 94470 47796
rect 100662 47744 100668 47796
rect 100720 47784 100726 47796
rect 106458 47784 106464 47796
rect 100720 47756 106464 47784
rect 100720 47744 100726 47756
rect 106458 47744 106464 47756
rect 106516 47744 106522 47796
rect 113082 47744 113088 47796
rect 113140 47784 113146 47796
rect 118510 47784 118516 47796
rect 113140 47756 118516 47784
rect 113140 47744 113146 47756
rect 118510 47744 118516 47756
rect 118568 47744 118574 47796
rect 121362 47744 121368 47796
rect 121420 47784 121426 47796
rect 126146 47784 126152 47796
rect 121420 47756 126152 47784
rect 121420 47744 121426 47756
rect 126146 47744 126152 47756
rect 126204 47744 126210 47796
rect 126882 47744 126888 47796
rect 126940 47784 126946 47796
rect 130562 47784 130568 47796
rect 126940 47756 130568 47784
rect 126940 47744 126946 47756
rect 130562 47744 130568 47756
rect 130620 47744 130626 47796
rect 132402 47744 132408 47796
rect 132460 47784 132466 47796
rect 135990 47784 135996 47796
rect 132460 47756 135996 47784
rect 132460 47744 132466 47756
rect 135990 47744 135996 47756
rect 136048 47744 136054 47796
rect 136542 47744 136548 47796
rect 136600 47784 136606 47796
rect 139302 47784 139308 47796
rect 136600 47756 139308 47784
rect 136600 47744 136606 47756
rect 139302 47744 139308 47756
rect 139360 47744 139366 47796
rect 147582 47744 147588 47796
rect 147640 47784 147646 47796
rect 150250 47784 150256 47796
rect 147640 47756 150256 47784
rect 147640 47744 147646 47756
rect 150250 47744 150256 47756
rect 150308 47744 150314 47796
rect 153010 47744 153016 47796
rect 153068 47784 153074 47796
rect 155678 47784 155684 47796
rect 153068 47756 155684 47784
rect 153068 47744 153074 47756
rect 155678 47744 155684 47756
rect 155736 47744 155742 47796
rect 193306 47744 193312 47796
rect 193364 47784 193370 47796
rect 194042 47784 194048 47796
rect 193364 47756 194048 47784
rect 193364 47744 193370 47756
rect 194042 47744 194048 47756
rect 194100 47744 194106 47796
rect 211614 47744 211620 47796
rect 211672 47784 211678 47796
rect 212718 47784 212724 47796
rect 211672 47756 212724 47784
rect 211672 47744 211678 47756
rect 212718 47744 212724 47756
rect 212776 47744 212782 47796
rect 225782 47744 225788 47796
rect 225840 47784 225846 47796
rect 227806 47784 227812 47796
rect 225840 47756 227812 47784
rect 225840 47744 225846 47756
rect 227806 47744 227812 47756
rect 227864 47744 227870 47796
rect 243354 47744 243360 47796
rect 243412 47784 243418 47796
rect 246298 47784 246304 47796
rect 243412 47756 246304 47784
rect 243412 47744 243418 47756
rect 246298 47744 246304 47756
rect 246356 47744 246362 47796
rect 306926 47744 306932 47796
rect 306984 47784 306990 47796
rect 307662 47784 307668 47796
rect 306984 47756 307668 47784
rect 306984 47744 306990 47756
rect 307662 47744 307668 47756
rect 307720 47744 307726 47796
rect 318978 47744 318984 47796
rect 319036 47784 319042 47796
rect 320082 47784 320088 47796
rect 319036 47756 320088 47784
rect 319036 47744 319042 47756
rect 320082 47744 320088 47756
rect 320140 47744 320146 47796
rect 370406 47744 370412 47796
rect 370464 47784 370470 47796
rect 371142 47784 371148 47796
rect 370464 47756 371148 47784
rect 370464 47744 370470 47756
rect 371142 47744 371148 47756
rect 371200 47744 371206 47796
rect 435082 47744 435088 47796
rect 435140 47784 435146 47796
rect 436002 47784 436008 47796
rect 435140 47756 436008 47784
rect 435140 47744 435146 47756
rect 436002 47744 436008 47756
rect 436060 47744 436066 47796
rect 534718 47744 534724 47796
rect 534776 47784 534782 47796
rect 536944 47784 536972 47824
rect 560938 47812 560944 47824
rect 560996 47812 561002 47864
rect 534776 47756 536972 47784
rect 534776 47744 534782 47756
rect 538030 47744 538036 47796
rect 538088 47784 538094 47796
rect 564526 47784 564532 47796
rect 538088 47756 564532 47784
rect 538088 47744 538094 47756
rect 564526 47744 564532 47756
rect 564584 47744 564590 47796
rect 66220 47688 74534 47716
rect 66220 47676 66226 47688
rect 85482 47676 85488 47728
rect 85540 47716 85546 47728
rect 92198 47716 92204 47728
rect 85540 47688 92204 47716
rect 85540 47676 85546 47688
rect 92198 47676 92204 47688
rect 92256 47676 92262 47728
rect 103422 47676 103428 47728
rect 103480 47716 103486 47728
rect 109678 47716 109684 47728
rect 103480 47688 109684 47716
rect 103480 47676 103486 47688
rect 109678 47676 109684 47688
rect 109736 47676 109742 47728
rect 111610 47676 111616 47728
rect 111668 47716 111674 47728
rect 116302 47716 116308 47728
rect 111668 47688 116308 47716
rect 111668 47676 111674 47688
rect 116302 47676 116308 47688
rect 116360 47676 116366 47728
rect 117222 47676 117228 47728
rect 117280 47716 117286 47728
rect 121730 47716 121736 47728
rect 117280 47688 121736 47716
rect 117280 47676 117286 47688
rect 121730 47676 121736 47688
rect 121788 47676 121794 47728
rect 122742 47676 122748 47728
rect 122800 47716 122806 47728
rect 127250 47716 127256 47728
rect 122800 47688 127256 47716
rect 122800 47676 122806 47688
rect 127250 47676 127256 47688
rect 127308 47676 127314 47728
rect 137922 47676 137928 47728
rect 137980 47716 137986 47728
rect 141510 47716 141516 47728
rect 137980 47688 141516 47716
rect 137980 47676 137986 47688
rect 141510 47676 141516 47688
rect 141568 47676 141574 47728
rect 238938 47676 238944 47728
rect 238996 47716 239002 47728
rect 240042 47716 240048 47728
rect 238996 47688 240048 47716
rect 238996 47676 239002 47688
rect 240042 47676 240048 47688
rect 240100 47676 240106 47728
rect 340874 47676 340880 47728
rect 340932 47716 340938 47728
rect 342070 47716 342076 47728
rect 340932 47688 342076 47716
rect 340932 47676 340938 47688
rect 342070 47676 342076 47688
rect 342128 47676 342134 47728
rect 498562 47676 498568 47728
rect 498620 47716 498626 47728
rect 502978 47716 502984 47728
rect 498620 47688 502984 47716
rect 498620 47676 498626 47688
rect 502978 47676 502984 47688
rect 503036 47676 503042 47728
rect 509510 47676 509516 47728
rect 509568 47716 509574 47728
rect 510522 47716 510528 47728
rect 509568 47688 510528 47716
rect 509568 47676 509574 47688
rect 510522 47676 510528 47688
rect 510580 47676 510586 47728
rect 528186 47676 528192 47728
rect 528244 47716 528250 47728
rect 549993 47719 550051 47725
rect 549993 47716 550005 47719
rect 528244 47688 550005 47716
rect 528244 47676 528250 47688
rect 549993 47685 550005 47688
rect 550039 47685 550051 47719
rect 549993 47679 550051 47685
rect 552290 47676 552296 47728
rect 552348 47716 552354 47728
rect 553302 47716 553308 47728
rect 552348 47688 553308 47716
rect 552348 47676 552354 47688
rect 553302 47676 553308 47688
rect 553360 47676 553366 47728
rect 66088 47620 69336 47648
rect 1302 47540 1308 47592
rect 1360 47580 1366 47592
rect 14458 47580 14464 47592
rect 1360 47552 14464 47580
rect 1360 47540 1366 47552
rect 14458 47540 14464 47552
rect 14516 47540 14522 47592
rect 20530 47540 20536 47592
rect 20588 47580 20594 47592
rect 32766 47580 32772 47592
rect 20588 47552 32772 47580
rect 20588 47540 20594 47552
rect 32766 47540 32772 47552
rect 32824 47540 32830 47592
rect 37182 47540 37188 47592
rect 37240 47580 37246 47592
rect 48406 47580 48412 47592
rect 37240 47552 48412 47580
rect 37240 47540 37246 47552
rect 48406 47540 48412 47552
rect 48464 47540 48470 47592
rect 49602 47540 49608 47592
rect 49660 47580 49666 47592
rect 59354 47580 59360 47592
rect 49660 47552 59360 47580
rect 49660 47540 49666 47552
rect 59354 47540 59360 47552
rect 59412 47540 59418 47592
rect 60642 47540 60648 47592
rect 60700 47580 60706 47592
rect 69198 47580 69204 47592
rect 60700 47552 69204 47580
rect 60700 47540 60706 47552
rect 69198 47540 69204 47552
rect 69256 47540 69262 47592
rect 10962 47472 10968 47524
rect 11020 47512 11026 47524
rect 23198 47512 23204 47524
rect 11020 47484 23204 47512
rect 11020 47472 11026 47484
rect 23198 47472 23204 47484
rect 23256 47472 23262 47524
rect 34422 47472 34428 47524
rect 34480 47512 34486 47524
rect 45094 47512 45100 47524
rect 34480 47484 45100 47512
rect 34480 47472 34486 47484
rect 45094 47472 45100 47484
rect 45152 47472 45158 47524
rect 69308 47512 69336 47620
rect 71682 47608 71688 47660
rect 71740 47648 71746 47660
rect 80146 47648 80152 47660
rect 71740 47620 80152 47648
rect 71740 47608 71746 47620
rect 80146 47608 80152 47620
rect 80204 47608 80210 47660
rect 81342 47608 81348 47660
rect 81400 47648 81406 47660
rect 88886 47648 88892 47660
rect 81400 47620 88892 47648
rect 81400 47608 81406 47620
rect 88886 47608 88892 47620
rect 88944 47608 88950 47660
rect 89622 47608 89628 47660
rect 89680 47648 89686 47660
rect 96614 47648 96620 47660
rect 89680 47620 96620 47648
rect 89680 47608 89686 47620
rect 96614 47608 96620 47620
rect 96672 47608 96678 47660
rect 104802 47608 104808 47660
rect 104860 47648 104866 47660
rect 110782 47648 110788 47660
rect 104860 47620 110788 47648
rect 104860 47608 104866 47620
rect 110782 47608 110788 47620
rect 110840 47608 110846 47660
rect 111702 47608 111708 47660
rect 111760 47648 111766 47660
rect 117406 47648 117412 47660
rect 111760 47620 117412 47648
rect 111760 47608 111766 47620
rect 117406 47608 117412 47620
rect 117464 47608 117470 47660
rect 157242 47608 157248 47660
rect 157300 47648 157306 47660
rect 158990 47648 158996 47660
rect 157300 47620 158996 47648
rect 157300 47608 157306 47620
rect 158990 47608 158996 47620
rect 159048 47608 159054 47660
rect 164142 47608 164148 47660
rect 164200 47648 164206 47660
rect 165614 47648 165620 47660
rect 164200 47620 165620 47648
rect 164200 47608 164206 47620
rect 165614 47608 165620 47620
rect 165672 47608 165678 47660
rect 218146 47608 218152 47660
rect 218204 47648 218210 47660
rect 219342 47648 219348 47660
rect 218204 47620 219348 47648
rect 218204 47608 218210 47620
rect 219342 47608 219348 47620
rect 219400 47608 219406 47660
rect 221458 47608 221464 47660
rect 221516 47648 221522 47660
rect 222838 47648 222844 47660
rect 221516 47620 222844 47648
rect 221516 47608 221522 47620
rect 222838 47608 222844 47620
rect 222896 47608 222902 47660
rect 223666 47608 223672 47660
rect 223724 47648 223730 47660
rect 224770 47648 224776 47660
rect 223724 47620 224776 47648
rect 223724 47608 223730 47620
rect 224770 47608 224776 47620
rect 224828 47608 224834 47660
rect 266354 47608 266360 47660
rect 266412 47648 266418 47660
rect 267642 47648 267648 47660
rect 266412 47620 267648 47648
rect 266412 47608 266418 47620
rect 267642 47608 267648 47620
rect 267700 47608 267706 47660
rect 276198 47608 276204 47660
rect 276256 47648 276262 47660
rect 277302 47648 277308 47660
rect 276256 47620 277308 47648
rect 276256 47608 276262 47620
rect 277302 47608 277308 47620
rect 277360 47608 277366 47660
rect 313458 47608 313464 47660
rect 313516 47648 313522 47660
rect 314562 47648 314568 47660
rect 313516 47620 314568 47648
rect 313516 47608 313522 47620
rect 314562 47608 314568 47620
rect 314620 47608 314626 47660
rect 356146 47608 356152 47660
rect 356204 47648 356210 47660
rect 357342 47648 357348 47660
rect 356204 47620 357348 47648
rect 356204 47608 356210 47620
rect 357342 47608 357348 47620
rect 357400 47608 357406 47660
rect 361666 47608 361672 47660
rect 361724 47648 361730 47660
rect 362862 47648 362868 47660
rect 361724 47620 362868 47648
rect 361724 47608 361730 47620
rect 362862 47608 362868 47620
rect 362920 47608 362926 47660
rect 495250 47608 495256 47660
rect 495308 47648 495314 47660
rect 504358 47648 504364 47660
rect 495308 47620 504364 47648
rect 495308 47608 495314 47620
rect 504358 47608 504364 47620
rect 504416 47608 504422 47660
rect 505186 47608 505192 47660
rect 505244 47648 505250 47660
rect 515398 47648 515404 47660
rect 505244 47620 515404 47648
rect 505244 47608 505250 47620
rect 515398 47608 515404 47620
rect 515456 47608 515462 47660
rect 541342 47608 541348 47660
rect 541400 47648 541406 47660
rect 568574 47648 568580 47660
rect 541400 47620 568580 47648
rect 541400 47608 541406 47620
rect 568574 47608 568580 47620
rect 568632 47608 568638 47660
rect 70210 47540 70216 47592
rect 70268 47580 70274 47592
rect 79042 47580 79048 47592
rect 70268 47552 79048 47580
rect 70268 47540 70274 47552
rect 79042 47540 79048 47552
rect 79100 47540 79106 47592
rect 82722 47540 82728 47592
rect 82780 47580 82786 47592
rect 89990 47580 89996 47592
rect 82780 47552 89996 47580
rect 82780 47540 82786 47552
rect 89990 47540 89996 47552
rect 90048 47540 90054 47592
rect 106182 47540 106188 47592
rect 106240 47580 106246 47592
rect 111886 47580 111892 47592
rect 106240 47552 111892 47580
rect 106240 47540 106246 47552
rect 111886 47540 111892 47552
rect 111944 47540 111950 47592
rect 259822 47540 259828 47592
rect 259880 47580 259886 47592
rect 260742 47580 260748 47592
rect 259880 47552 260748 47580
rect 259880 47540 259886 47552
rect 260742 47540 260748 47552
rect 260800 47540 260806 47592
rect 265250 47540 265256 47592
rect 265308 47580 265314 47592
rect 270586 47580 270592 47592
rect 265308 47552 270592 47580
rect 265308 47540 265314 47552
rect 270586 47540 270592 47552
rect 270644 47540 270650 47592
rect 275094 47540 275100 47592
rect 275152 47580 275158 47592
rect 275922 47580 275928 47592
rect 275152 47552 275928 47580
rect 275152 47540 275158 47552
rect 275922 47540 275928 47552
rect 275980 47540 275986 47592
rect 280614 47540 280620 47592
rect 280672 47580 280678 47592
rect 281442 47580 281448 47592
rect 280672 47552 281448 47580
rect 280672 47540 280678 47552
rect 281442 47540 281448 47552
rect 281500 47540 281506 47592
rect 323302 47540 323308 47592
rect 323360 47580 323366 47592
rect 324222 47580 324228 47592
rect 323360 47552 324228 47580
rect 323360 47540 323366 47552
rect 324222 47540 324228 47552
rect 324280 47540 324286 47592
rect 344094 47540 344100 47592
rect 344152 47580 344158 47592
rect 344922 47580 344928 47592
rect 344152 47552 344928 47580
rect 344152 47540 344158 47552
rect 344922 47540 344928 47552
rect 344980 47540 344986 47592
rect 349614 47540 349620 47592
rect 349672 47580 349678 47592
rect 350442 47580 350448 47592
rect 349672 47552 350448 47580
rect 349672 47540 349678 47552
rect 350442 47540 350448 47552
rect 350500 47540 350506 47592
rect 381354 47540 381360 47592
rect 381412 47580 381418 47592
rect 382182 47580 382188 47592
rect 381412 47552 382188 47580
rect 381412 47540 381418 47552
rect 382182 47540 382188 47552
rect 382240 47540 382246 47592
rect 397822 47540 397828 47592
rect 397880 47580 397886 47592
rect 398742 47580 398748 47592
rect 397880 47552 398748 47580
rect 397880 47540 397886 47552
rect 398742 47540 398748 47552
rect 398800 47540 398806 47592
rect 424134 47540 424140 47592
rect 424192 47580 424198 47592
rect 424962 47580 424968 47592
rect 424192 47552 424968 47580
rect 424192 47540 424198 47552
rect 424962 47540 424968 47552
rect 425020 47540 425026 47592
rect 444926 47540 444932 47592
rect 444984 47580 444990 47592
rect 445662 47580 445668 47592
rect 444984 47552 445668 47580
rect 444984 47540 444990 47552
rect 445662 47540 445668 47552
rect 445720 47540 445726 47592
rect 455874 47540 455880 47592
rect 455932 47580 455938 47592
rect 456702 47580 456708 47592
rect 455932 47552 456708 47580
rect 455932 47540 455938 47552
rect 456702 47540 456708 47552
rect 456760 47540 456766 47592
rect 462406 47540 462412 47592
rect 462464 47580 462470 47592
rect 482278 47580 482284 47592
rect 462464 47552 482284 47580
rect 462464 47540 462470 47552
rect 482278 47540 482284 47552
rect 482336 47540 482342 47592
rect 487614 47540 487620 47592
rect 487672 47580 487678 47592
rect 488442 47580 488448 47592
rect 487672 47552 488448 47580
rect 487672 47540 487678 47552
rect 488442 47540 488448 47552
rect 488500 47540 488506 47592
rect 488718 47540 488724 47592
rect 488776 47580 488782 47592
rect 512086 47580 512092 47592
rect 488776 47552 512092 47580
rect 488776 47540 488782 47552
rect 512086 47540 512092 47552
rect 512144 47540 512150 47592
rect 553394 47540 553400 47592
rect 553452 47580 553458 47592
rect 582377 47583 582435 47589
rect 582377 47580 582389 47583
rect 553452 47552 582389 47580
rect 553452 47540 553458 47552
rect 582377 47549 582389 47552
rect 582423 47549 582435 47583
rect 582377 47543 582435 47549
rect 73522 47512 73528 47524
rect 69308 47484 73528 47512
rect 73522 47472 73528 47484
rect 73580 47472 73586 47524
rect 393406 47472 393412 47524
rect 393464 47512 393470 47524
rect 394510 47512 394516 47524
rect 393464 47484 394516 47512
rect 393464 47472 393470 47484
rect 394510 47472 394516 47484
rect 394568 47472 394574 47524
rect 549993 47515 550051 47521
rect 549993 47481 550005 47515
rect 550039 47512 550051 47515
rect 554774 47512 554780 47524
rect 550039 47484 554780 47512
rect 550039 47481 550051 47484
rect 549993 47475 550051 47481
rect 554774 47472 554780 47484
rect 554832 47472 554838 47524
rect 15102 47404 15108 47456
rect 15160 47444 15166 47456
rect 27522 47444 27528 47456
rect 15160 47416 27528 47444
rect 15160 47404 15166 47416
rect 27522 47404 27528 47416
rect 27580 47404 27586 47456
rect 75822 47404 75828 47456
rect 75880 47444 75886 47456
rect 83458 47444 83464 47456
rect 75880 47416 83464 47444
rect 75880 47404 75886 47416
rect 83458 47404 83464 47416
rect 83516 47404 83522 47456
rect 96522 47404 96528 47456
rect 96580 47444 96586 47456
rect 103146 47444 103152 47456
rect 96580 47416 103152 47444
rect 96580 47404 96586 47416
rect 103146 47404 103152 47416
rect 103204 47404 103210 47456
rect 143442 47404 143448 47456
rect 143500 47444 143506 47456
rect 145834 47444 145840 47456
rect 143500 47416 145840 47444
rect 143500 47404 143506 47416
rect 145834 47404 145840 47416
rect 145892 47404 145898 47456
rect 345198 47404 345204 47456
rect 345256 47444 345262 47456
rect 346302 47444 346308 47456
rect 345256 47416 346308 47444
rect 345256 47404 345262 47416
rect 346302 47404 346308 47416
rect 346360 47404 346366 47456
rect 398926 47404 398932 47456
rect 398984 47444 398990 47456
rect 400030 47444 400036 47456
rect 398984 47416 400036 47444
rect 398984 47404 398990 47416
rect 400030 47404 400036 47416
rect 400088 47404 400094 47456
rect 414198 47404 414204 47456
rect 414256 47444 414262 47456
rect 415302 47444 415308 47456
rect 414256 47416 415308 47444
rect 414256 47404 414262 47416
rect 415302 47404 415308 47416
rect 415360 47404 415366 47456
rect 425238 47404 425244 47456
rect 425296 47444 425302 47456
rect 426342 47444 426348 47456
rect 425296 47416 426348 47444
rect 425296 47404 425302 47416
rect 426342 47404 426348 47416
rect 426400 47404 426406 47456
rect 447134 47404 447140 47456
rect 447192 47444 447198 47456
rect 448422 47444 448428 47456
rect 447192 47416 448428 47444
rect 447192 47404 447198 47416
rect 448422 47404 448428 47416
rect 448480 47404 448486 47456
rect 16482 47336 16488 47388
rect 16540 47376 16546 47388
rect 28626 47376 28632 47388
rect 16540 47348 28632 47376
rect 16540 47336 16546 47348
rect 28626 47336 28632 47348
rect 28684 47336 28690 47388
rect 22002 47268 22008 47320
rect 22060 47308 22066 47320
rect 34146 47308 34152 47320
rect 22060 47280 34152 47308
rect 22060 47268 22066 47280
rect 34146 47268 34152 47280
rect 34204 47268 34210 47320
rect 95142 47268 95148 47320
rect 95200 47308 95206 47320
rect 100938 47308 100944 47320
rect 95200 47280 100944 47308
rect 95200 47268 95206 47280
rect 100938 47268 100944 47280
rect 100996 47268 101002 47320
rect 124122 47268 124128 47320
rect 124180 47308 124186 47320
rect 128354 47308 128360 47320
rect 124180 47280 128360 47308
rect 124180 47268 124186 47280
rect 128354 47268 128360 47280
rect 128412 47268 128418 47320
rect 207198 47268 207204 47320
rect 207256 47308 207262 47320
rect 208486 47308 208492 47320
rect 207256 47280 208492 47308
rect 207256 47268 207262 47280
rect 208486 47268 208492 47280
rect 208544 47268 208550 47320
rect 298094 47268 298100 47320
rect 298152 47308 298158 47320
rect 299290 47308 299296 47320
rect 298152 47280 299296 47308
rect 298152 47268 298158 47280
rect 299290 47268 299296 47280
rect 299348 47268 299354 47320
rect 492030 47268 492036 47320
rect 492088 47308 492094 47320
rect 497458 47308 497464 47320
rect 492088 47280 497464 47308
rect 492088 47268 492094 47280
rect 497458 47268 497464 47280
rect 497516 47268 497522 47320
rect 542446 47268 542452 47320
rect 542504 47308 542510 47320
rect 543642 47308 543648 47320
rect 542504 47280 543648 47308
rect 542504 47268 542510 47280
rect 543642 47268 543648 47280
rect 543700 47268 543706 47320
rect 119890 47132 119896 47184
rect 119948 47172 119954 47184
rect 125042 47172 125048 47184
rect 119948 47144 125048 47172
rect 119948 47132 119954 47144
rect 125042 47132 125048 47144
rect 125100 47132 125106 47184
rect 128262 47132 128268 47184
rect 128320 47172 128326 47184
rect 132678 47172 132684 47184
rect 128320 47144 132684 47172
rect 128320 47132 128326 47144
rect 132678 47132 132684 47144
rect 132736 47132 132742 47184
rect 110322 47064 110328 47116
rect 110380 47104 110386 47116
rect 115198 47104 115204 47116
rect 110380 47076 115204 47104
rect 110380 47064 110386 47076
rect 115198 47064 115204 47076
rect 115256 47064 115262 47116
rect 131022 47064 131028 47116
rect 131080 47104 131086 47116
rect 134886 47104 134892 47116
rect 131080 47076 134892 47104
rect 131080 47064 131086 47076
rect 134886 47064 134892 47076
rect 134944 47064 134950 47116
rect 139302 47064 139308 47116
rect 139360 47104 139366 47116
rect 142614 47104 142620 47116
rect 139360 47076 142620 47104
rect 139360 47064 139366 47076
rect 142614 47064 142620 47076
rect 142672 47064 142678 47116
rect 78490 46996 78496 47048
rect 78548 47036 78554 47048
rect 86678 47036 86684 47048
rect 78548 47008 86684 47036
rect 78548 46996 78554 47008
rect 86678 46996 86684 47008
rect 86736 46996 86742 47048
rect 99282 46996 99288 47048
rect 99340 47036 99346 47048
rect 105354 47036 105360 47048
rect 99340 47008 105360 47036
rect 99340 46996 99346 47008
rect 105354 46996 105360 47008
rect 105412 46996 105418 47048
rect 108942 46996 108948 47048
rect 109000 47036 109006 47048
rect 114094 47036 114100 47048
rect 109000 47008 114100 47036
rect 109000 46996 109006 47008
rect 114094 46996 114100 47008
rect 114152 46996 114158 47048
rect 118602 46996 118608 47048
rect 118660 47036 118666 47048
rect 122834 47036 122840 47048
rect 118660 47008 122840 47036
rect 118660 46996 118666 47008
rect 122834 46996 122840 47008
rect 122892 46996 122898 47048
rect 125502 46996 125508 47048
rect 125560 47036 125566 47048
rect 129458 47036 129464 47048
rect 125560 47008 129464 47036
rect 125560 46996 125566 47008
rect 129458 46996 129464 47008
rect 129516 46996 129522 47048
rect 129642 46996 129648 47048
rect 129700 47036 129706 47048
rect 133782 47036 133788 47048
rect 129700 47008 133788 47036
rect 129700 46996 129706 47008
rect 133782 46996 133788 47008
rect 133840 46996 133846 47048
rect 140682 46996 140688 47048
rect 140740 47036 140746 47048
rect 143626 47036 143632 47048
rect 140740 47008 143632 47036
rect 140740 46996 140746 47008
rect 143626 46996 143632 47008
rect 143684 46996 143690 47048
rect 151722 46996 151728 47048
rect 151780 47036 151786 47048
rect 153562 47036 153568 47048
rect 151780 47008 153568 47036
rect 151780 46996 151786 47008
rect 153562 46996 153568 47008
rect 153620 46996 153626 47048
rect 271874 46996 271880 47048
rect 271932 47036 271938 47048
rect 277486 47036 277492 47048
rect 271932 47008 277492 47036
rect 271932 46996 271938 47008
rect 277486 46996 277492 47008
rect 277544 46996 277550 47048
rect 68922 46928 68928 46980
rect 68980 46968 68986 46980
rect 76834 46968 76840 46980
rect 68980 46940 76840 46968
rect 68980 46928 68986 46940
rect 76834 46928 76840 46940
rect 76892 46928 76898 46980
rect 78582 46928 78588 46980
rect 78640 46968 78646 46980
rect 85574 46968 85580 46980
rect 78640 46940 85580 46968
rect 78640 46928 78646 46940
rect 85574 46928 85580 46940
rect 85632 46928 85638 46980
rect 88242 46928 88248 46980
rect 88300 46968 88306 46980
rect 95510 46968 95516 46980
rect 88300 46940 95516 46968
rect 88300 46928 88306 46940
rect 95510 46928 95516 46940
rect 95568 46928 95574 46980
rect 97902 46928 97908 46980
rect 97960 46968 97966 46980
rect 104250 46968 104256 46980
rect 97960 46940 104256 46968
rect 97960 46928 97966 46940
rect 104250 46928 104256 46940
rect 104308 46928 104314 46980
rect 119982 46928 119988 46980
rect 120040 46968 120046 46980
rect 123938 46968 123944 46980
rect 120040 46940 123944 46968
rect 120040 46928 120046 46940
rect 123938 46928 123944 46940
rect 123996 46928 124002 46980
rect 137094 46968 137100 46980
rect 133800 46940 137100 46968
rect 133800 46912 133828 46940
rect 137094 46928 137100 46940
rect 137152 46928 137158 46980
rect 142062 46928 142068 46980
rect 142120 46968 142126 46980
rect 144730 46968 144736 46980
rect 142120 46940 144736 46968
rect 142120 46928 142126 46940
rect 144730 46928 144736 46940
rect 144788 46928 144794 46980
rect 148042 46968 148048 46980
rect 144840 46940 148048 46968
rect 133782 46860 133788 46912
rect 133840 46860 133846 46912
rect 144840 46776 144868 46940
rect 148042 46928 148048 46940
rect 148100 46928 148106 46980
rect 151078 46928 151084 46980
rect 151136 46968 151142 46980
rect 152458 46968 152464 46980
rect 151136 46940 152464 46968
rect 151136 46928 151142 46940
rect 152458 46928 152464 46940
rect 152516 46928 152522 46980
rect 161290 46928 161296 46980
rect 161348 46968 161354 46980
rect 163406 46968 163412 46980
rect 161348 46940 163412 46968
rect 161348 46928 161354 46940
rect 163406 46928 163412 46940
rect 163464 46928 163470 46980
rect 199562 46928 199568 46980
rect 199620 46968 199626 46980
rect 200206 46968 200212 46980
rect 199620 46940 200212 46968
rect 199620 46928 199626 46940
rect 200206 46928 200212 46940
rect 200264 46928 200270 46980
rect 219250 46928 219256 46980
rect 219308 46968 219314 46980
rect 220078 46968 220084 46980
rect 219308 46940 220084 46968
rect 219308 46928 219314 46940
rect 220078 46928 220084 46940
rect 220136 46928 220142 46980
rect 566458 46860 566464 46912
rect 566516 46900 566522 46912
rect 580166 46900 580172 46912
rect 566516 46872 580172 46900
rect 566516 46860 566522 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 144822 46724 144828 46776
rect 144880 46724 144886 46776
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 7558 45540 7564 45552
rect 3568 45512 7564 45540
rect 3568 45500 3574 45512
rect 7558 45500 7564 45512
rect 7616 45500 7622 45552
rect 558178 33056 558184 33108
rect 558236 33096 558242 33108
rect 580166 33096 580172 33108
rect 558236 33068 580172 33096
rect 558236 33056 558242 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 2774 32920 2780 32972
rect 2832 32960 2838 32972
rect 6178 32960 6184 32972
rect 2832 32932 6184 32960
rect 2832 32920 2838 32932
rect 6178 32920 6184 32932
rect 6236 32920 6242 32972
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 10318 20652 10324 20664
rect 3568 20624 10324 20652
rect 3568 20612 3574 20624
rect 10318 20612 10324 20624
rect 10376 20612 10382 20664
rect 562318 20612 562324 20664
rect 562376 20652 562382 20664
rect 579982 20652 579988 20664
rect 562376 20624 579988 20652
rect 562376 20612 562382 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 474550 11840 474556 11892
rect 474608 11840 474614 11892
rect 474568 11676 474596 11840
rect 474642 11676 474648 11688
rect 474568 11648 474648 11676
rect 474642 11636 474648 11648
rect 474700 11636 474706 11688
rect 515398 7692 515404 7744
rect 515456 7732 515462 7744
rect 530118 7732 530124 7744
rect 515456 7704 530124 7732
rect 515456 7692 515462 7704
rect 530118 7692 530124 7704
rect 530176 7692 530182 7744
rect 480070 7624 480076 7676
rect 480128 7664 480134 7676
rect 501782 7664 501788 7676
rect 480128 7636 501788 7664
rect 480128 7624 480134 7636
rect 501782 7624 501788 7636
rect 501840 7624 501846 7676
rect 504358 7624 504364 7676
rect 504416 7664 504422 7676
rect 519538 7664 519544 7676
rect 504416 7636 519544 7664
rect 504416 7624 504422 7636
rect 519538 7624 519544 7636
rect 519596 7624 519602 7676
rect 469030 7556 469036 7608
rect 469088 7596 469094 7608
rect 491110 7596 491116 7608
rect 469088 7568 491116 7596
rect 469088 7556 469094 7568
rect 491110 7556 491116 7568
rect 491168 7556 491174 7608
rect 497458 7556 497464 7608
rect 497516 7596 497522 7608
rect 515950 7596 515956 7608
rect 497516 7568 515956 7596
rect 497516 7556 497522 7568
rect 515950 7556 515956 7568
rect 516008 7556 516014 7608
rect 516042 7556 516048 7608
rect 516100 7596 516106 7608
rect 540790 7596 540796 7608
rect 516100 7568 540796 7596
rect 516100 7556 516106 7568
rect 540790 7556 540796 7568
rect 540848 7556 540854 7608
rect 556798 6808 556804 6860
rect 556856 6848 556862 6860
rect 580166 6848 580172 6860
rect 556856 6820 580172 6848
rect 556856 6808 556862 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 560938 5516 560944 5568
rect 560996 5556 561002 5568
rect 562042 5556 562048 5568
rect 560996 5528 562048 5556
rect 560996 5516 561002 5528
rect 562042 5516 562048 5528
rect 562100 5516 562106 5568
rect 502978 5176 502984 5228
rect 503036 5216 503042 5228
rect 523034 5216 523040 5228
rect 503036 5188 523040 5216
rect 503036 5176 503042 5188
rect 523034 5176 523040 5188
rect 523092 5176 523098 5228
rect 509142 5108 509148 5160
rect 509200 5148 509206 5160
rect 533706 5148 533712 5160
rect 509200 5120 533712 5148
rect 509200 5108 509206 5120
rect 533706 5108 533712 5120
rect 533764 5108 533770 5160
rect 473262 5040 473268 5092
rect 473320 5080 473326 5092
rect 494698 5080 494704 5092
rect 473320 5052 494704 5080
rect 473320 5040 473326 5052
rect 494698 5040 494704 5052
rect 494756 5040 494762 5092
rect 502242 5040 502248 5092
rect 502300 5080 502306 5092
rect 526622 5080 526628 5092
rect 502300 5052 526628 5080
rect 502300 5040 502306 5052
rect 526622 5040 526628 5052
rect 526680 5040 526686 5092
rect 466362 4972 466368 5024
rect 466420 5012 466426 5024
rect 487614 5012 487620 5024
rect 466420 4984 487620 5012
rect 466420 4972 466426 4984
rect 487614 4972 487620 4984
rect 487672 4972 487678 5024
rect 518802 4972 518808 5024
rect 518860 5012 518866 5024
rect 544378 5012 544384 5024
rect 518860 4984 544384 5012
rect 518860 4972 518866 4984
rect 544378 4972 544384 4984
rect 544436 4972 544442 5024
rect 485682 4904 485688 4956
rect 485740 4944 485746 4956
rect 508866 4944 508872 4956
rect 485740 4916 508872 4944
rect 485740 4904 485746 4916
rect 508866 4904 508872 4916
rect 508924 4904 508930 4956
rect 525702 4904 525708 4956
rect 525760 4944 525766 4956
rect 551462 4944 551468 4956
rect 525760 4916 551468 4944
rect 525760 4904 525766 4916
rect 551462 4904 551468 4916
rect 551520 4904 551526 4956
rect 476022 4836 476028 4888
rect 476080 4876 476086 4888
rect 498194 4876 498200 4888
rect 476080 4848 498200 4876
rect 476080 4836 476086 4848
rect 498194 4836 498200 4848
rect 498252 4836 498258 4888
rect 511810 4836 511816 4888
rect 511868 4876 511874 4888
rect 537202 4876 537208 4888
rect 511868 4848 537208 4876
rect 511868 4836 511874 4848
rect 537202 4836 537208 4848
rect 537260 4836 537266 4888
rect 459462 4768 459468 4820
rect 459520 4808 459526 4820
rect 480530 4808 480536 4820
rect 459520 4780 480536 4808
rect 459520 4768 459526 4780
rect 480530 4768 480536 4780
rect 480588 4768 480594 4820
rect 482922 4768 482928 4820
rect 482980 4808 482986 4820
rect 505370 4808 505376 4820
rect 482980 4780 505376 4808
rect 482980 4768 482986 4780
rect 505370 4768 505376 4780
rect 505428 4768 505434 4820
rect 521470 4768 521476 4820
rect 521528 4808 521534 4820
rect 547874 4808 547880 4820
rect 521528 4780 547880 4808
rect 521528 4768 521534 4780
rect 547874 4768 547880 4780
rect 547932 4768 547938 4820
rect 482278 4156 482284 4208
rect 482336 4196 482342 4208
rect 484026 4196 484032 4208
rect 482336 4168 484032 4196
rect 482336 4156 482342 4168
rect 484026 4156 484032 4168
rect 484084 4156 484090 4208
rect 209682 4088 209688 4140
rect 209740 4128 209746 4140
rect 210970 4128 210976 4140
rect 209740 4100 210976 4128
rect 209740 4088 209746 4100
rect 210970 4088 210976 4100
rect 211028 4088 211034 4140
rect 229002 4088 229008 4140
rect 229060 4128 229066 4140
rect 231026 4128 231032 4140
rect 229060 4100 231032 4128
rect 229060 4088 229066 4100
rect 231026 4088 231032 4100
rect 231084 4088 231090 4140
rect 237282 4088 237288 4140
rect 237340 4128 237346 4140
rect 240502 4128 240508 4140
rect 237340 4100 240508 4128
rect 237340 4088 237346 4100
rect 240502 4088 240508 4100
rect 240560 4088 240566 4140
rect 256510 4088 256516 4140
rect 256568 4128 256574 4140
rect 260650 4128 260656 4140
rect 256568 4100 260656 4128
rect 256568 4088 256574 4100
rect 260650 4088 260656 4100
rect 260708 4088 260714 4140
rect 262122 4088 262128 4140
rect 262180 4128 262186 4140
rect 267734 4128 267740 4140
rect 262180 4100 267740 4128
rect 262180 4088 262186 4100
rect 267734 4088 267740 4100
rect 267792 4088 267798 4140
rect 282730 4088 282736 4140
rect 282788 4128 282794 4140
rect 288986 4128 288992 4140
rect 282788 4100 288992 4128
rect 282788 4088 282794 4100
rect 288986 4088 288992 4100
rect 289044 4088 289050 4140
rect 323302 4128 323308 4140
rect 316006 4100 323308 4128
rect 253842 4020 253848 4072
rect 253900 4060 253906 4072
rect 258258 4060 258264 4072
rect 253900 4032 258264 4060
rect 253900 4020 253906 4032
rect 258258 4020 258264 4032
rect 258316 4020 258322 4072
rect 304902 4020 304908 4072
rect 304960 4060 304966 4072
rect 312630 4060 312636 4072
rect 304960 4032 312636 4060
rect 304960 4020 304966 4032
rect 312630 4020 312636 4032
rect 312688 4020 312694 4072
rect 314562 4020 314568 4072
rect 314620 4060 314626 4072
rect 316006 4060 316034 4100
rect 323302 4088 323308 4100
rect 323360 4088 323366 4140
rect 324222 4088 324228 4140
rect 324280 4128 324286 4140
rect 333882 4128 333888 4140
rect 324280 4100 333888 4128
rect 324280 4088 324286 4100
rect 333882 4088 333888 4100
rect 333940 4088 333946 4140
rect 343542 4088 343548 4140
rect 343600 4128 343606 4140
rect 355226 4128 355232 4140
rect 343600 4100 355232 4128
rect 343600 4088 343606 4100
rect 355226 4088 355232 4100
rect 355284 4088 355290 4140
rect 355962 4088 355968 4140
rect 356020 4128 356026 4140
rect 368198 4128 368204 4140
rect 356020 4100 368204 4128
rect 356020 4088 356026 4100
rect 368198 4088 368204 4100
rect 368256 4088 368262 4140
rect 371142 4088 371148 4140
rect 371200 4128 371206 4140
rect 384758 4128 384764 4140
rect 371200 4100 384764 4128
rect 371200 4088 371206 4100
rect 384758 4088 384764 4100
rect 384816 4088 384822 4140
rect 384942 4088 384948 4140
rect 385000 4128 385006 4140
rect 399938 4128 399944 4140
rect 385000 4100 399944 4128
rect 385000 4088 385006 4100
rect 399938 4088 399944 4100
rect 399996 4088 400002 4140
rect 411070 4088 411076 4140
rect 411128 4128 411134 4140
rect 427262 4128 427268 4140
rect 411128 4100 427268 4128
rect 411128 4088 411134 4100
rect 427262 4088 427268 4100
rect 427320 4088 427326 4140
rect 429102 4088 429108 4140
rect 429160 4128 429166 4140
rect 447410 4128 447416 4140
rect 429160 4100 447416 4128
rect 429160 4088 429166 4100
rect 447410 4088 447416 4100
rect 447468 4088 447474 4140
rect 451182 4088 451188 4140
rect 451240 4128 451246 4140
rect 471054 4128 471060 4140
rect 451240 4100 471060 4128
rect 451240 4088 451246 4100
rect 471054 4088 471060 4100
rect 471112 4088 471118 4140
rect 477402 4088 477408 4140
rect 477460 4128 477466 4140
rect 499390 4128 499396 4140
rect 477460 4100 499396 4128
rect 477460 4088 477466 4100
rect 499390 4088 499396 4100
rect 499448 4088 499454 4140
rect 505002 4088 505008 4140
rect 505060 4128 505066 4140
rect 529014 4128 529020 4140
rect 505060 4100 529020 4128
rect 505060 4088 505066 4100
rect 529014 4088 529020 4100
rect 529072 4088 529078 4140
rect 529842 4088 529848 4140
rect 529900 4128 529906 4140
rect 556154 4128 556160 4140
rect 529900 4100 556160 4128
rect 529900 4088 529906 4100
rect 556154 4088 556160 4100
rect 556212 4088 556218 4140
rect 320910 4060 320916 4072
rect 314620 4032 316034 4060
rect 317248 4032 320916 4060
rect 314620 4020 314626 4032
rect 245470 3952 245476 4004
rect 245528 3992 245534 4004
rect 249978 3992 249984 4004
rect 245528 3964 249984 3992
rect 245528 3952 245534 3964
rect 249978 3952 249984 3964
rect 250036 3952 250042 4004
rect 264882 3952 264888 4004
rect 264940 3992 264946 4004
rect 270034 3992 270040 4004
rect 264940 3964 270040 3992
rect 264940 3952 264946 3964
rect 270034 3952 270040 3964
rect 270092 3952 270098 4004
rect 281442 3952 281448 4004
rect 281500 3992 281506 4004
rect 287790 3992 287796 4004
rect 281500 3964 287796 3992
rect 281500 3952 281506 3964
rect 287790 3952 287796 3964
rect 287848 3952 287854 4004
rect 293770 3952 293776 4004
rect 293828 3992 293834 4004
rect 300762 3992 300768 4004
rect 293828 3964 300768 3992
rect 293828 3952 293834 3964
rect 300762 3952 300768 3964
rect 300820 3952 300826 4004
rect 311802 3952 311808 4004
rect 311860 3992 311866 4004
rect 317248 3992 317276 4032
rect 320910 4020 320916 4032
rect 320968 4020 320974 4072
rect 331122 4020 331128 4072
rect 331180 4060 331186 4072
rect 340966 4060 340972 4072
rect 331180 4032 340972 4060
rect 331180 4020 331186 4032
rect 340966 4020 340972 4032
rect 341024 4020 341030 4072
rect 342070 4020 342076 4072
rect 342128 4060 342134 4072
rect 352834 4060 352840 4072
rect 342128 4032 352840 4060
rect 342128 4020 342134 4032
rect 352834 4020 352840 4032
rect 352892 4020 352898 4072
rect 354582 4020 354588 4072
rect 354640 4060 354646 4072
rect 366910 4060 366916 4072
rect 354640 4032 366916 4060
rect 354640 4020 354646 4032
rect 366910 4020 366916 4032
rect 366968 4020 366974 4072
rect 373810 4020 373816 4072
rect 373868 4060 373874 4072
rect 387150 4060 387156 4072
rect 373868 4032 387156 4060
rect 373868 4020 373874 4032
rect 387150 4020 387156 4032
rect 387208 4020 387214 4072
rect 394510 4020 394516 4072
rect 394568 4060 394574 4072
rect 409598 4060 409604 4072
rect 394568 4032 409604 4060
rect 394568 4020 394574 4032
rect 409598 4020 409604 4032
rect 409656 4020 409662 4072
rect 416682 4020 416688 4072
rect 416740 4060 416746 4072
rect 434438 4060 434444 4072
rect 416740 4032 434444 4060
rect 416740 4020 416746 4032
rect 434438 4020 434444 4032
rect 434496 4020 434502 4072
rect 434622 4020 434628 4072
rect 434680 4060 434686 4072
rect 453298 4060 453304 4072
rect 434680 4032 453304 4060
rect 434680 4020 434686 4032
rect 453298 4020 453304 4032
rect 453356 4020 453362 4072
rect 456702 4020 456708 4072
rect 456760 4060 456766 4072
rect 476942 4060 476948 4072
rect 456760 4032 476948 4060
rect 456760 4020 456766 4032
rect 476942 4020 476948 4032
rect 477000 4020 477006 4072
rect 481542 4020 481548 4072
rect 481600 4060 481606 4072
rect 504174 4060 504180 4072
rect 481600 4032 504180 4060
rect 481600 4020 481606 4032
rect 504174 4020 504180 4032
rect 504232 4020 504238 4072
rect 510522 4020 510528 4072
rect 510580 4060 510586 4072
rect 534902 4060 534908 4072
rect 510580 4032 534908 4060
rect 510580 4020 510586 4032
rect 534902 4020 534908 4032
rect 534960 4020 534966 4072
rect 543642 4020 543648 4072
rect 543700 4060 543706 4072
rect 570322 4060 570328 4072
rect 543700 4032 570328 4060
rect 543700 4020 543706 4032
rect 570322 4020 570328 4032
rect 570380 4020 570386 4072
rect 311860 3964 317276 3992
rect 311860 3952 311866 3964
rect 317322 3952 317328 4004
rect 317380 3952 317386 4004
rect 332502 3952 332508 4004
rect 332560 3992 332566 4004
rect 343358 3992 343364 4004
rect 332560 3964 343364 3992
rect 332560 3952 332566 3964
rect 343358 3952 343364 3964
rect 343416 3952 343422 4004
rect 346302 3952 346308 4004
rect 346360 3992 346366 4004
rect 357526 3992 357532 4004
rect 346360 3964 357532 3992
rect 346360 3952 346366 3964
rect 357526 3952 357532 3964
rect 357584 3952 357590 4004
rect 365622 3952 365628 4004
rect 365680 3992 365686 4004
rect 378870 3992 378876 4004
rect 365680 3964 378876 3992
rect 365680 3952 365686 3964
rect 378870 3952 378876 3964
rect 378928 3952 378934 4004
rect 382182 3952 382188 4004
rect 382240 3992 382246 4004
rect 396534 3992 396540 4004
rect 382240 3964 396540 3992
rect 382240 3952 382246 3964
rect 396534 3952 396540 3964
rect 396592 3952 396598 4004
rect 398742 3952 398748 4004
rect 398800 3992 398806 4004
rect 414290 3992 414296 4004
rect 398800 3964 414296 3992
rect 398800 3952 398806 3964
rect 414290 3952 414296 3964
rect 414348 3952 414354 4004
rect 420730 3952 420736 4004
rect 420788 3992 420794 4004
rect 437934 3992 437940 4004
rect 420788 3964 437940 3992
rect 420788 3952 420794 3964
rect 437934 3952 437940 3964
rect 437992 3952 437998 4004
rect 441522 3952 441528 4004
rect 441580 3992 441586 4004
rect 460382 3992 460388 4004
rect 441580 3964 460388 3992
rect 441580 3952 441586 3964
rect 460382 3952 460388 3964
rect 460440 3952 460446 4004
rect 463602 3952 463608 4004
rect 463660 3992 463666 4004
rect 485222 3992 485228 4004
rect 463660 3964 485228 3992
rect 463660 3952 463666 3964
rect 485222 3952 485228 3964
rect 485280 3952 485286 4004
rect 487062 3952 487068 4004
rect 487120 3992 487126 4004
rect 510062 3992 510068 4004
rect 487120 3964 510068 3992
rect 487120 3952 487126 3964
rect 510062 3952 510068 3964
rect 510120 3952 510126 4004
rect 514662 3952 514668 4004
rect 514720 3992 514726 4004
rect 539594 3992 539600 4004
rect 514720 3964 539600 3992
rect 514720 3952 514726 3964
rect 539594 3952 539600 3964
rect 539652 3952 539658 4004
rect 546402 3952 546408 4004
rect 546460 3992 546466 4004
rect 573910 3992 573916 4004
rect 546460 3964 573916 3992
rect 546460 3952 546466 3964
rect 573910 3952 573916 3964
rect 573968 3952 573974 4004
rect 303522 3884 303528 3936
rect 303580 3924 303586 3936
rect 311434 3924 311440 3936
rect 303580 3896 311440 3924
rect 303580 3884 303586 3896
rect 311434 3884 311440 3896
rect 311492 3884 311498 3936
rect 317340 3924 317368 3952
rect 326798 3924 326804 3936
rect 317340 3896 326804 3924
rect 326798 3884 326804 3896
rect 326856 3884 326862 3936
rect 326982 3884 326988 3936
rect 327040 3924 327046 3936
rect 337470 3924 337476 3936
rect 327040 3896 337476 3924
rect 327040 3884 327046 3896
rect 337470 3884 337476 3896
rect 337528 3884 337534 3936
rect 342162 3884 342168 3936
rect 342220 3924 342226 3936
rect 354030 3924 354036 3936
rect 342220 3896 354036 3924
rect 342220 3884 342226 3896
rect 354030 3884 354036 3896
rect 354088 3884 354094 3936
rect 354646 3896 360056 3924
rect 248322 3816 248328 3868
rect 248380 3856 248386 3868
rect 252370 3856 252376 3868
rect 248380 3828 252376 3856
rect 248380 3816 248386 3828
rect 252370 3816 252376 3828
rect 252428 3816 252434 3868
rect 274542 3816 274548 3868
rect 274600 3856 274606 3868
rect 280706 3856 280712 3868
rect 274600 3828 280712 3856
rect 274600 3816 274606 3828
rect 280706 3816 280712 3828
rect 280764 3816 280770 3868
rect 292482 3816 292488 3868
rect 292540 3856 292546 3868
rect 299658 3856 299664 3868
rect 292540 3828 299664 3856
rect 292540 3816 292546 3828
rect 299658 3816 299664 3828
rect 299716 3816 299722 3868
rect 308950 3816 308956 3868
rect 309008 3856 309014 3868
rect 317322 3856 317328 3868
rect 309008 3828 317328 3856
rect 309008 3816 309014 3828
rect 317322 3816 317328 3828
rect 317380 3816 317386 3868
rect 318702 3816 318708 3868
rect 318760 3856 318766 3868
rect 327994 3856 328000 3868
rect 318760 3828 328000 3856
rect 318760 3816 318766 3828
rect 327994 3816 328000 3828
rect 328052 3816 328058 3868
rect 328362 3816 328368 3868
rect 328420 3856 328426 3868
rect 338666 3856 338672 3868
rect 328420 3828 338672 3856
rect 328420 3816 328426 3828
rect 338666 3816 338672 3828
rect 338724 3816 338730 3868
rect 339402 3816 339408 3868
rect 339460 3856 339466 3868
rect 350442 3856 350448 3868
rect 339460 3828 350448 3856
rect 339460 3816 339466 3828
rect 350442 3816 350448 3828
rect 350500 3816 350506 3868
rect 351730 3816 351736 3868
rect 351788 3856 351794 3868
rect 354646 3856 354674 3896
rect 359918 3856 359924 3868
rect 351788 3828 354674 3856
rect 358648 3828 359924 3856
rect 351788 3816 351794 3828
rect 286962 3748 286968 3800
rect 287020 3788 287026 3800
rect 293678 3788 293684 3800
rect 287020 3760 293684 3788
rect 287020 3748 287026 3760
rect 293678 3748 293684 3760
rect 293736 3748 293742 3800
rect 309042 3748 309048 3800
rect 309100 3788 309106 3800
rect 318518 3788 318524 3800
rect 309100 3760 318524 3788
rect 309100 3748 309106 3760
rect 318518 3748 318524 3760
rect 318576 3748 318582 3800
rect 320082 3748 320088 3800
rect 320140 3788 320146 3800
rect 329190 3788 329196 3800
rect 320140 3760 329196 3788
rect 320140 3748 320146 3760
rect 329190 3748 329196 3760
rect 329248 3748 329254 3800
rect 329742 3748 329748 3800
rect 329800 3788 329806 3800
rect 339862 3788 339868 3800
rect 329800 3760 339868 3788
rect 329800 3748 329806 3760
rect 339862 3748 339868 3760
rect 339920 3748 339926 3800
rect 347682 3748 347688 3800
rect 347740 3788 347746 3800
rect 358648 3788 358676 3828
rect 359918 3816 359924 3828
rect 359976 3816 359982 3868
rect 360028 3856 360056 3896
rect 360102 3884 360108 3936
rect 360160 3924 360166 3936
rect 372890 3924 372896 3936
rect 360160 3896 372896 3924
rect 360160 3884 360166 3896
rect 372890 3884 372896 3896
rect 372948 3884 372954 3936
rect 373902 3884 373908 3936
rect 373960 3924 373966 3936
rect 388254 3924 388260 3936
rect 373960 3896 388260 3924
rect 373960 3884 373966 3896
rect 388254 3884 388260 3896
rect 388312 3884 388318 3936
rect 394602 3884 394608 3936
rect 394660 3924 394666 3936
rect 410794 3924 410800 3936
rect 394660 3896 410800 3924
rect 394660 3884 394666 3896
rect 410794 3884 410800 3896
rect 410852 3884 410858 3936
rect 412542 3884 412548 3936
rect 412600 3924 412606 3936
rect 429654 3924 429660 3936
rect 412600 3896 429660 3924
rect 412600 3884 412606 3896
rect 429654 3884 429660 3896
rect 429712 3884 429718 3936
rect 430482 3884 430488 3936
rect 430540 3924 430546 3936
rect 448606 3924 448612 3936
rect 430540 3896 448612 3924
rect 430540 3884 430546 3896
rect 448606 3884 448612 3896
rect 448664 3884 448670 3936
rect 457990 3884 457996 3936
rect 458048 3924 458054 3936
rect 478138 3924 478144 3936
rect 458048 3896 478144 3924
rect 458048 3884 458054 3896
rect 478138 3884 478144 3896
rect 478196 3884 478202 3936
rect 484302 3884 484308 3936
rect 484360 3924 484366 3936
rect 507670 3924 507676 3936
rect 484360 3896 507676 3924
rect 484360 3884 484366 3896
rect 507670 3884 507676 3896
rect 507728 3884 507734 3936
rect 507762 3884 507768 3936
rect 507820 3924 507826 3936
rect 532510 3924 532516 3936
rect 507820 3896 532516 3924
rect 507820 3884 507826 3896
rect 532510 3884 532516 3896
rect 532568 3884 532574 3936
rect 539502 3884 539508 3936
rect 539560 3924 539566 3936
rect 566826 3924 566832 3936
rect 539560 3896 566832 3924
rect 539560 3884 539566 3896
rect 566826 3884 566832 3896
rect 566884 3884 566890 3936
rect 363506 3856 363512 3868
rect 360028 3828 363512 3856
rect 363506 3816 363512 3828
rect 363564 3816 363570 3868
rect 367002 3816 367008 3868
rect 367060 3856 367066 3868
rect 379974 3856 379980 3868
rect 367060 3828 379980 3856
rect 367060 3816 367066 3828
rect 379974 3816 379980 3828
rect 380032 3816 380038 3868
rect 383470 3816 383476 3868
rect 383528 3856 383534 3868
rect 397730 3856 397736 3868
rect 383528 3828 397736 3856
rect 383528 3816 383534 3828
rect 397730 3816 397736 3828
rect 397788 3816 397794 3868
rect 400122 3816 400128 3868
rect 400180 3856 400186 3868
rect 416682 3856 416688 3868
rect 400180 3828 416688 3856
rect 400180 3816 400186 3828
rect 416682 3816 416688 3828
rect 416740 3816 416746 3868
rect 422202 3816 422208 3868
rect 422260 3856 422266 3868
rect 440326 3856 440332 3868
rect 422260 3828 440332 3856
rect 422260 3816 422266 3828
rect 440326 3816 440332 3828
rect 440384 3816 440390 3868
rect 444282 3816 444288 3868
rect 444340 3856 444346 3868
rect 463970 3856 463976 3868
rect 444340 3828 463976 3856
rect 444340 3816 444346 3828
rect 463970 3816 463976 3828
rect 464028 3816 464034 3868
rect 470502 3816 470508 3868
rect 470560 3856 470566 3868
rect 492306 3856 492312 3868
rect 470560 3828 492312 3856
rect 470560 3816 470566 3828
rect 492306 3816 492312 3828
rect 492364 3816 492370 3868
rect 493962 3816 493968 3868
rect 494020 3856 494026 3868
rect 517146 3856 517152 3868
rect 494020 3828 517152 3856
rect 494020 3816 494026 3828
rect 517146 3816 517152 3828
rect 517204 3816 517210 3868
rect 521562 3816 521568 3868
rect 521620 3856 521626 3868
rect 546678 3856 546684 3868
rect 521620 3828 546684 3856
rect 521620 3816 521626 3828
rect 546678 3816 546684 3828
rect 546736 3816 546742 3868
rect 549070 3816 549076 3868
rect 549128 3856 549134 3868
rect 576302 3856 576308 3868
rect 549128 3828 576308 3856
rect 549128 3816 549134 3828
rect 576302 3816 576308 3828
rect 576360 3816 576366 3868
rect 347740 3760 358676 3788
rect 347740 3748 347746 3760
rect 358722 3748 358728 3800
rect 358780 3788 358786 3800
rect 358780 3760 358860 3788
rect 358780 3748 358786 3760
rect 235902 3680 235908 3732
rect 235960 3720 235966 3732
rect 239306 3720 239312 3732
rect 235960 3692 239312 3720
rect 235960 3680 235966 3692
rect 239306 3680 239312 3692
rect 239364 3680 239370 3732
rect 267642 3680 267648 3732
rect 267700 3720 267706 3732
rect 272426 3720 272432 3732
rect 267700 3692 272432 3720
rect 267700 3680 267706 3692
rect 272426 3680 272432 3692
rect 272484 3680 272490 3732
rect 275922 3680 275928 3732
rect 275980 3720 275986 3732
rect 281902 3720 281908 3732
rect 275980 3692 281908 3720
rect 275980 3680 275986 3692
rect 281902 3680 281908 3692
rect 281960 3680 281966 3732
rect 284202 3680 284208 3732
rect 284260 3720 284266 3732
rect 291378 3720 291384 3732
rect 284260 3692 291384 3720
rect 284260 3680 284266 3692
rect 291378 3680 291384 3692
rect 291436 3680 291442 3732
rect 295242 3680 295248 3732
rect 295300 3720 295306 3732
rect 303154 3720 303160 3732
rect 295300 3692 303160 3720
rect 295300 3680 295306 3692
rect 303154 3680 303160 3692
rect 303212 3680 303218 3732
rect 306282 3680 306288 3732
rect 306340 3720 306346 3732
rect 315022 3720 315028 3732
rect 306340 3692 315028 3720
rect 306340 3680 306346 3692
rect 315022 3680 315028 3692
rect 315080 3680 315086 3732
rect 315942 3680 315948 3732
rect 316000 3720 316006 3732
rect 316000 3692 325464 3720
rect 316000 3680 316006 3692
rect 238662 3612 238668 3664
rect 238720 3652 238726 3664
rect 241698 3652 241704 3664
rect 238720 3624 241704 3652
rect 238720 3612 238726 3624
rect 241698 3612 241704 3624
rect 241756 3612 241762 3664
rect 257982 3612 257988 3664
rect 258040 3652 258046 3664
rect 262950 3652 262956 3664
rect 258040 3624 262956 3652
rect 258040 3612 258046 3624
rect 262950 3612 262956 3624
rect 263008 3612 263014 3664
rect 277302 3612 277308 3664
rect 277360 3652 277366 3664
rect 283098 3652 283104 3664
rect 277360 3624 283104 3652
rect 277360 3612 277366 3624
rect 283098 3612 283104 3624
rect 283156 3612 283162 3664
rect 285582 3612 285588 3664
rect 285640 3652 285646 3664
rect 292574 3652 292580 3664
rect 285640 3624 292580 3652
rect 285640 3612 285646 3624
rect 292574 3612 292580 3624
rect 292632 3612 292638 3664
rect 293862 3612 293868 3664
rect 293920 3652 293926 3664
rect 301958 3652 301964 3664
rect 293920 3624 301964 3652
rect 293920 3612 293926 3624
rect 301958 3612 301964 3624
rect 302016 3612 302022 3664
rect 302142 3612 302148 3664
rect 302200 3652 302206 3664
rect 310238 3652 310244 3664
rect 302200 3624 310244 3652
rect 302200 3612 302206 3624
rect 310238 3612 310244 3624
rect 310296 3612 310302 3664
rect 313182 3612 313188 3664
rect 313240 3652 313246 3664
rect 322106 3652 322112 3664
rect 313240 3624 322112 3652
rect 313240 3612 313246 3624
rect 322106 3612 322112 3624
rect 322164 3612 322170 3664
rect 325436 3652 325464 3692
rect 325510 3680 325516 3732
rect 325568 3720 325574 3732
rect 335078 3720 335084 3732
rect 325568 3692 335084 3720
rect 325568 3680 325574 3692
rect 335078 3680 335084 3692
rect 335136 3680 335142 3732
rect 336642 3680 336648 3732
rect 336700 3720 336706 3732
rect 346946 3720 346952 3732
rect 336700 3692 346952 3720
rect 336700 3680 336706 3692
rect 346946 3680 346952 3692
rect 347004 3680 347010 3732
rect 349062 3680 349068 3732
rect 349120 3720 349126 3732
rect 358633 3723 358691 3729
rect 358633 3720 358645 3723
rect 349120 3692 358645 3720
rect 349120 3680 349126 3692
rect 358633 3689 358645 3692
rect 358679 3689 358691 3723
rect 358633 3683 358691 3689
rect 325602 3652 325608 3664
rect 325436 3624 325608 3652
rect 325602 3612 325608 3624
rect 325660 3612 325666 3664
rect 331030 3612 331036 3664
rect 331088 3652 331094 3664
rect 331088 3624 332824 3652
rect 331088 3612 331094 3624
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 3970 3584 3976 3596
rect 2924 3556 3976 3584
rect 2924 3544 2930 3556
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 20530 3584 20536 3596
rect 19484 3556 20536 3584
rect 19484 3544 19490 3556
rect 20530 3544 20536 3556
rect 20588 3544 20594 3596
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 28810 3584 28816 3596
rect 27764 3556 28816 3584
rect 27764 3544 27770 3556
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45370 3584 45376 3596
rect 44324 3556 45376 3584
rect 44324 3544 44330 3556
rect 45370 3544 45376 3556
rect 45428 3544 45434 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 70210 3584 70216 3596
rect 69164 3556 70216 3584
rect 69164 3544 69170 3556
rect 70210 3544 70216 3556
rect 70268 3544 70274 3596
rect 77386 3544 77392 3596
rect 77444 3584 77450 3596
rect 78490 3584 78496 3596
rect 77444 3556 78496 3584
rect 77444 3544 77450 3556
rect 78490 3544 78496 3556
rect 78548 3544 78554 3596
rect 93946 3544 93952 3596
rect 94004 3584 94010 3596
rect 95050 3584 95056 3596
rect 94004 3556 95056 3584
rect 94004 3544 94010 3556
rect 95050 3544 95056 3556
rect 95108 3544 95114 3596
rect 168374 3544 168380 3596
rect 168432 3584 168438 3596
rect 169662 3584 169668 3596
rect 168432 3556 169668 3584
rect 168432 3544 168438 3556
rect 169662 3544 169668 3556
rect 169720 3544 169726 3596
rect 186314 3544 186320 3596
rect 186372 3584 186378 3596
rect 187326 3584 187332 3596
rect 186372 3556 187332 3584
rect 186372 3544 186378 3556
rect 187326 3544 187332 3556
rect 187384 3544 187390 3596
rect 201494 3544 201500 3596
rect 201552 3584 201558 3596
rect 202690 3584 202696 3596
rect 201552 3556 202696 3584
rect 201552 3544 201558 3556
rect 202690 3544 202696 3556
rect 202748 3544 202754 3596
rect 219342 3544 219348 3596
rect 219400 3584 219406 3596
rect 220446 3584 220452 3596
rect 219400 3556 220452 3584
rect 219400 3544 219406 3556
rect 220446 3544 220452 3556
rect 220504 3544 220510 3596
rect 223482 3544 223488 3596
rect 223540 3584 223546 3596
rect 225138 3584 225144 3596
rect 223540 3556 225144 3584
rect 223540 3544 223546 3556
rect 225138 3544 225144 3556
rect 225196 3544 225202 3596
rect 242802 3544 242808 3596
rect 242860 3584 242866 3596
rect 246390 3584 246396 3596
rect 242860 3556 246396 3584
rect 242860 3544 242866 3556
rect 246390 3544 246396 3556
rect 246448 3544 246454 3596
rect 251082 3544 251088 3596
rect 251140 3584 251146 3596
rect 255866 3584 255872 3596
rect 251140 3556 255872 3584
rect 251140 3544 251146 3556
rect 255866 3544 255872 3556
rect 255924 3544 255930 3596
rect 282822 3544 282828 3596
rect 282880 3584 282886 3596
rect 290182 3584 290188 3596
rect 282880 3556 290188 3584
rect 282880 3544 282886 3556
rect 290182 3544 290188 3556
rect 290240 3544 290246 3596
rect 299382 3544 299388 3596
rect 299440 3584 299446 3596
rect 307938 3584 307944 3596
rect 299440 3556 307944 3584
rect 299440 3544 299446 3556
rect 307938 3544 307944 3556
rect 307996 3544 308002 3596
rect 310422 3544 310428 3596
rect 310480 3584 310486 3596
rect 319714 3584 319720 3596
rect 310480 3556 319720 3584
rect 310480 3544 310486 3556
rect 319714 3544 319720 3556
rect 319772 3544 319778 3596
rect 322842 3544 322848 3596
rect 322900 3584 322906 3596
rect 332686 3584 332692 3596
rect 322900 3556 332692 3584
rect 322900 3544 322906 3556
rect 332686 3544 332692 3556
rect 332744 3544 332750 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12250 3516 12256 3528
rect 11204 3488 12256 3516
rect 11204 3476 11210 3488
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 37090 3516 37096 3528
rect 36044 3488 37096 3516
rect 36044 3476 36050 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 52362 3516 52368 3528
rect 51408 3488 52368 3516
rect 51408 3476 51414 3488
rect 52362 3476 52368 3488
rect 52420 3476 52426 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 53650 3516 53656 3528
rect 52604 3488 53656 3516
rect 52604 3476 52610 3488
rect 53650 3476 53656 3488
rect 53708 3476 53714 3528
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 56502 3516 56508 3528
rect 56100 3488 56508 3516
rect 56100 3476 56106 3488
rect 56502 3476 56508 3488
rect 56560 3476 56566 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 60826 3476 60832 3528
rect 60884 3516 60890 3528
rect 61930 3516 61936 3528
rect 60884 3488 61936 3516
rect 60884 3476 60890 3488
rect 61930 3476 61936 3488
rect 61988 3476 61994 3528
rect 64322 3476 64328 3528
rect 64380 3516 64386 3528
rect 64782 3516 64788 3528
rect 64380 3488 64788 3516
rect 64380 3476 64386 3488
rect 64782 3476 64788 3488
rect 64840 3476 64846 3528
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 66714 3476 66720 3528
rect 66772 3516 66778 3528
rect 67542 3516 67548 3528
rect 66772 3488 67548 3516
rect 66772 3476 66778 3488
rect 67542 3476 67548 3488
rect 67600 3476 67606 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 82078 3476 82084 3528
rect 82136 3516 82142 3528
rect 82722 3516 82728 3528
rect 82136 3488 82728 3516
rect 82136 3476 82142 3488
rect 82722 3476 82728 3488
rect 82780 3476 82786 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 92382 3516 92388 3528
rect 91612 3488 92388 3516
rect 91612 3476 91618 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 102042 3516 102048 3528
rect 101088 3488 102048 3516
rect 101088 3476 101094 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 102226 3476 102232 3528
rect 102284 3516 102290 3528
rect 103238 3516 103244 3528
rect 102284 3488 103244 3516
rect 102284 3476 102290 3488
rect 103238 3476 103244 3488
rect 103296 3476 103302 3528
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 106182 3516 106188 3528
rect 105780 3488 106188 3516
rect 105780 3476 105786 3488
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 110322 3516 110328 3528
rect 109368 3488 110328 3516
rect 109368 3476 109374 3488
rect 110322 3476 110328 3488
rect 110380 3476 110386 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111518 3516 111524 3528
rect 110564 3488 111524 3516
rect 110564 3476 110570 3488
rect 111518 3476 111524 3488
rect 111576 3476 111582 3528
rect 114002 3476 114008 3528
rect 114060 3516 114066 3528
rect 114462 3516 114468 3528
rect 114060 3488 114468 3516
rect 114060 3476 114066 3488
rect 114462 3476 114468 3488
rect 114520 3476 114526 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 116394 3476 116400 3528
rect 116452 3516 116458 3528
rect 117222 3516 117228 3528
rect 116452 3488 117228 3516
rect 116452 3476 116458 3488
rect 117222 3476 117228 3488
rect 117280 3476 117286 3528
rect 117590 3476 117596 3528
rect 117648 3516 117654 3528
rect 118602 3516 118608 3528
rect 117648 3488 118608 3516
rect 117648 3476 117654 3488
rect 118602 3476 118608 3488
rect 118660 3476 118666 3528
rect 118786 3476 118792 3528
rect 118844 3516 118850 3528
rect 119982 3516 119988 3528
rect 118844 3488 119988 3516
rect 118844 3476 118850 3488
rect 119982 3476 119988 3488
rect 120040 3476 120046 3528
rect 122282 3476 122288 3528
rect 122340 3516 122346 3528
rect 122742 3516 122748 3528
rect 122340 3488 122748 3516
rect 122340 3476 122346 3488
rect 122742 3476 122748 3488
rect 122800 3476 122806 3528
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 126882 3516 126888 3528
rect 125928 3488 126888 3516
rect 125928 3476 125934 3488
rect 126882 3476 126888 3488
rect 126940 3476 126946 3528
rect 130562 3476 130568 3528
rect 130620 3516 130626 3528
rect 131022 3516 131028 3528
rect 130620 3488 131028 3516
rect 130620 3476 130626 3488
rect 131022 3476 131028 3488
rect 131080 3476 131086 3528
rect 132954 3476 132960 3528
rect 133012 3516 133018 3528
rect 133782 3516 133788 3528
rect 133012 3488 133788 3516
rect 133012 3476 133018 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
rect 134150 3476 134156 3528
rect 134208 3516 134214 3528
rect 135162 3516 135168 3528
rect 134208 3488 135168 3516
rect 134208 3476 134214 3488
rect 135162 3476 135168 3488
rect 135220 3476 135226 3528
rect 136450 3476 136456 3528
rect 136508 3516 136514 3528
rect 137278 3516 137284 3528
rect 136508 3488 137284 3516
rect 136508 3476 136514 3488
rect 137278 3476 137284 3488
rect 137336 3476 137342 3528
rect 138842 3476 138848 3528
rect 138900 3516 138906 3528
rect 139302 3516 139308 3528
rect 138900 3488 139308 3516
rect 138900 3476 138906 3488
rect 139302 3476 139308 3488
rect 139360 3476 139366 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 140682 3516 140688 3528
rect 140096 3488 140688 3516
rect 140096 3476 140102 3488
rect 140682 3476 140688 3488
rect 140740 3476 140746 3528
rect 141234 3476 141240 3528
rect 141292 3516 141298 3528
rect 142062 3516 142068 3528
rect 141292 3488 142068 3516
rect 141292 3476 141298 3488
rect 142062 3476 142068 3488
rect 142120 3476 142126 3528
rect 142430 3476 142436 3528
rect 142488 3516 142494 3528
rect 143442 3516 143448 3528
rect 142488 3488 143448 3516
rect 142488 3476 142494 3488
rect 143442 3476 143448 3488
rect 143500 3476 143506 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 148318 3476 148324 3528
rect 148376 3516 148382 3528
rect 148962 3516 148968 3528
rect 148376 3488 148968 3516
rect 148376 3476 148382 3488
rect 148962 3476 148968 3488
rect 149020 3476 149026 3528
rect 149514 3476 149520 3528
rect 149572 3516 149578 3528
rect 151078 3516 151084 3528
rect 149572 3488 151084 3516
rect 149572 3476 149578 3488
rect 151078 3476 151084 3488
rect 151136 3476 151142 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 153102 3516 153108 3528
rect 151872 3488 153108 3516
rect 151872 3476 151878 3488
rect 153102 3476 153108 3488
rect 153160 3476 153166 3528
rect 154206 3476 154212 3528
rect 154264 3516 154270 3528
rect 156046 3516 156052 3528
rect 154264 3488 156052 3516
rect 154264 3476 154270 3488
rect 156046 3476 156052 3488
rect 156104 3476 156110 3528
rect 156598 3476 156604 3528
rect 156656 3516 156662 3528
rect 157242 3516 157248 3528
rect 156656 3488 157248 3516
rect 156656 3476 156662 3488
rect 157242 3476 157248 3488
rect 157300 3476 157306 3528
rect 157794 3476 157800 3528
rect 157852 3516 157858 3528
rect 158622 3516 158628 3528
rect 157852 3488 158628 3516
rect 157852 3476 157858 3488
rect 158622 3476 158628 3488
rect 158680 3476 158686 3528
rect 158898 3476 158904 3528
rect 158956 3516 158962 3528
rect 160002 3516 160008 3528
rect 158956 3488 160008 3516
rect 158956 3476 158962 3488
rect 160002 3476 160008 3488
rect 160060 3476 160066 3528
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161382 3516 161388 3528
rect 160152 3488 161388 3516
rect 160152 3476 160158 3488
rect 161382 3476 161388 3488
rect 161440 3476 161446 3528
rect 163682 3476 163688 3528
rect 163740 3516 163746 3528
rect 164142 3516 164148 3528
rect 163740 3488 164148 3516
rect 163740 3476 163746 3488
rect 164142 3476 164148 3488
rect 164200 3476 164206 3528
rect 164878 3476 164884 3528
rect 164936 3516 164942 3528
rect 165706 3516 165712 3528
rect 164936 3488 165712 3516
rect 164936 3476 164942 3488
rect 165706 3476 165712 3488
rect 165764 3476 165770 3528
rect 166074 3476 166080 3528
rect 166132 3516 166138 3528
rect 166902 3516 166908 3528
rect 166132 3488 166908 3516
rect 166132 3476 166138 3488
rect 166902 3476 166908 3488
rect 166960 3476 166966 3528
rect 167178 3476 167184 3528
rect 167236 3516 167242 3528
rect 168558 3516 168564 3528
rect 167236 3488 168564 3516
rect 167236 3476 167242 3488
rect 168558 3476 168564 3488
rect 168616 3476 168622 3528
rect 171962 3476 171968 3528
rect 172020 3516 172026 3528
rect 172606 3516 172612 3528
rect 172020 3488 172612 3516
rect 172020 3476 172026 3488
rect 172606 3476 172612 3488
rect 172664 3476 172670 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173802 3516 173808 3528
rect 173216 3488 173808 3516
rect 173216 3476 173222 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 174262 3476 174268 3528
rect 174320 3516 174326 3528
rect 175182 3516 175188 3528
rect 174320 3488 175188 3516
rect 174320 3476 174326 3488
rect 175182 3476 175188 3488
rect 175240 3476 175246 3528
rect 179046 3476 179052 3528
rect 179104 3516 179110 3528
rect 179506 3516 179512 3528
rect 179104 3488 179512 3516
rect 179104 3476 179110 3488
rect 179506 3476 179512 3488
rect 179564 3476 179570 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180702 3516 180708 3528
rect 180300 3488 180708 3516
rect 180300 3476 180306 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 180978 3476 180984 3528
rect 181036 3516 181042 3528
rect 181438 3516 181444 3528
rect 181036 3488 181444 3516
rect 181036 3476 181042 3488
rect 181438 3476 181444 3488
rect 181496 3476 181502 3528
rect 187694 3476 187700 3528
rect 187752 3516 187758 3528
rect 188522 3516 188528 3528
rect 187752 3488 188528 3516
rect 187752 3476 187758 3488
rect 188522 3476 188528 3488
rect 188580 3476 188586 3528
rect 189074 3476 189080 3528
rect 189132 3516 189138 3528
rect 189718 3516 189724 3528
rect 189132 3488 189724 3516
rect 189132 3476 189138 3488
rect 189718 3476 189724 3488
rect 189776 3476 189782 3528
rect 194594 3476 194600 3528
rect 194652 3516 194658 3528
rect 195606 3516 195612 3528
rect 194652 3488 195612 3516
rect 194652 3476 194658 3488
rect 195606 3476 195612 3488
rect 195664 3476 195670 3528
rect 198642 3476 198648 3528
rect 198700 3516 198706 3528
rect 199102 3516 199108 3528
rect 198700 3488 199108 3516
rect 198700 3476 198706 3488
rect 199102 3476 199108 3488
rect 199160 3476 199166 3528
rect 202782 3476 202788 3528
rect 202840 3516 202846 3528
rect 203886 3516 203892 3528
rect 202840 3488 203892 3516
rect 202840 3476 202846 3488
rect 203886 3476 203892 3488
rect 203944 3476 203950 3528
rect 205542 3476 205548 3528
rect 205600 3516 205606 3528
rect 206186 3516 206192 3528
rect 205600 3488 206192 3516
rect 205600 3476 205606 3488
rect 206186 3476 206192 3488
rect 206244 3476 206250 3528
rect 206922 3476 206928 3528
rect 206980 3516 206986 3528
rect 207382 3516 207388 3528
rect 206980 3488 207388 3516
rect 206980 3476 206986 3488
rect 207382 3476 207388 3488
rect 207440 3476 207446 3528
rect 211062 3476 211068 3528
rect 211120 3516 211126 3528
rect 212166 3516 212172 3528
rect 211120 3488 212172 3516
rect 211120 3476 211126 3488
rect 212166 3476 212172 3488
rect 212224 3476 212230 3528
rect 215202 3476 215208 3528
rect 215260 3516 215266 3528
rect 216858 3516 216864 3528
rect 215260 3488 216864 3516
rect 215260 3476 215266 3488
rect 216858 3476 216864 3488
rect 216916 3476 216922 3528
rect 217962 3476 217968 3528
rect 218020 3516 218026 3528
rect 219250 3516 219256 3528
rect 218020 3488 219256 3516
rect 218020 3476 218026 3488
rect 219250 3476 219256 3488
rect 219308 3476 219314 3528
rect 220078 3476 220084 3528
rect 220136 3516 220142 3528
rect 221550 3516 221556 3528
rect 220136 3488 221556 3516
rect 220136 3476 220142 3488
rect 221550 3476 221556 3488
rect 221608 3476 221614 3528
rect 222838 3476 222844 3528
rect 222896 3516 222902 3528
rect 223942 3516 223948 3528
rect 222896 3488 223948 3516
rect 222896 3476 222902 3488
rect 223942 3476 223948 3488
rect 224000 3476 224006 3528
rect 227622 3476 227628 3528
rect 227680 3516 227686 3528
rect 229830 3516 229836 3528
rect 227680 3488 229836 3516
rect 227680 3476 227686 3488
rect 229830 3476 229836 3488
rect 229888 3476 229894 3528
rect 233142 3476 233148 3528
rect 233200 3516 233206 3528
rect 235810 3516 235816 3528
rect 233200 3488 235816 3516
rect 233200 3476 233206 3488
rect 235810 3476 235816 3488
rect 235868 3476 235874 3528
rect 240778 3476 240784 3528
rect 240836 3516 240842 3528
rect 244090 3516 244096 3528
rect 240836 3488 244096 3516
rect 240836 3476 240842 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 246942 3476 246948 3528
rect 247000 3516 247006 3528
rect 251174 3516 251180 3528
rect 247000 3488 251180 3516
rect 247000 3476 247006 3488
rect 251174 3476 251180 3488
rect 251232 3476 251238 3528
rect 256602 3476 256608 3528
rect 256660 3516 256666 3528
rect 261754 3516 261760 3528
rect 256660 3488 261760 3516
rect 256660 3476 256666 3488
rect 261754 3476 261760 3488
rect 261812 3476 261818 3528
rect 269022 3476 269028 3528
rect 269080 3516 269086 3528
rect 274818 3516 274824 3528
rect 269080 3488 274824 3516
rect 269080 3476 269086 3488
rect 274818 3476 274824 3488
rect 274876 3476 274882 3528
rect 289722 3476 289728 3528
rect 289780 3516 289786 3528
rect 297266 3516 297272 3528
rect 289780 3488 297272 3516
rect 289780 3476 289786 3488
rect 297266 3476 297272 3488
rect 297324 3476 297330 3528
rect 299290 3476 299296 3528
rect 299348 3516 299354 3528
rect 306742 3516 306748 3528
rect 299348 3488 306748 3516
rect 299348 3476 299354 3488
rect 306742 3476 306748 3488
rect 306800 3476 306806 3528
rect 307662 3476 307668 3528
rect 307720 3516 307726 3528
rect 316218 3516 316224 3528
rect 307720 3488 316224 3516
rect 307720 3476 307726 3488
rect 316218 3476 316224 3488
rect 316276 3476 316282 3528
rect 321462 3476 321468 3528
rect 321520 3516 321526 3528
rect 331582 3516 331588 3528
rect 321520 3488 331588 3516
rect 321520 3476 321526 3488
rect 331582 3476 331588 3488
rect 331640 3476 331646 3528
rect 332796 3516 332824 3624
rect 335262 3612 335268 3664
rect 335320 3652 335326 3664
rect 345750 3652 345756 3664
rect 335320 3624 345756 3652
rect 335320 3612 335326 3624
rect 345750 3612 345756 3624
rect 345808 3612 345814 3664
rect 346210 3612 346216 3664
rect 346268 3652 346274 3664
rect 358722 3652 358728 3664
rect 346268 3624 358728 3652
rect 346268 3612 346274 3624
rect 358722 3612 358728 3624
rect 358780 3612 358786 3664
rect 358832 3652 358860 3760
rect 361482 3748 361488 3800
rect 361540 3788 361546 3800
rect 374086 3788 374092 3800
rect 361540 3760 374092 3788
rect 361540 3748 361546 3760
rect 374086 3748 374092 3760
rect 374144 3748 374150 3800
rect 380802 3748 380808 3800
rect 380860 3788 380866 3800
rect 395338 3788 395344 3800
rect 380860 3760 395344 3788
rect 380860 3748 380866 3760
rect 395338 3748 395344 3760
rect 395396 3748 395402 3800
rect 395982 3748 395988 3800
rect 396040 3788 396046 3800
rect 411898 3788 411904 3800
rect 396040 3760 411904 3788
rect 396040 3748 396046 3760
rect 411898 3748 411904 3760
rect 411956 3748 411962 3800
rect 415302 3748 415308 3800
rect 415360 3788 415366 3800
rect 432046 3788 432052 3800
rect 415360 3760 432052 3788
rect 415360 3748 415366 3760
rect 432046 3748 432052 3760
rect 432104 3748 432110 3800
rect 437290 3748 437296 3800
rect 437348 3788 437354 3800
rect 455690 3788 455696 3800
rect 437348 3760 455696 3788
rect 437348 3748 437354 3760
rect 455690 3748 455696 3760
rect 455748 3748 455754 3800
rect 460842 3748 460848 3800
rect 460900 3788 460906 3800
rect 481726 3788 481732 3800
rect 460900 3760 481732 3788
rect 460900 3748 460906 3760
rect 481726 3748 481732 3760
rect 481784 3748 481790 3800
rect 484210 3748 484216 3800
rect 484268 3788 484274 3800
rect 506474 3788 506480 3800
rect 484268 3760 506480 3788
rect 484268 3748 484274 3760
rect 506474 3748 506480 3760
rect 506532 3748 506538 3800
rect 513282 3748 513288 3800
rect 513340 3788 513346 3800
rect 538398 3788 538404 3800
rect 513340 3760 538404 3788
rect 513340 3748 513346 3760
rect 538398 3748 538404 3760
rect 538456 3748 538462 3800
rect 545022 3748 545028 3800
rect 545080 3788 545086 3800
rect 572714 3788 572720 3800
rect 545080 3760 572720 3788
rect 545080 3748 545086 3760
rect 572714 3748 572720 3760
rect 572772 3748 572778 3800
rect 362770 3680 362776 3732
rect 362828 3720 362834 3732
rect 376478 3720 376484 3732
rect 362828 3692 376484 3720
rect 362828 3680 362834 3692
rect 376478 3680 376484 3692
rect 376536 3680 376542 3732
rect 376662 3680 376668 3732
rect 376720 3720 376726 3732
rect 390646 3720 390652 3732
rect 376720 3692 390652 3720
rect 376720 3680 376726 3692
rect 390646 3680 390652 3692
rect 390704 3680 390710 3732
rect 391842 3680 391848 3732
rect 391900 3720 391906 3732
rect 407206 3720 407212 3732
rect 391900 3692 407212 3720
rect 391900 3680 391906 3692
rect 407206 3680 407212 3692
rect 407264 3680 407270 3732
rect 411162 3680 411168 3732
rect 411220 3720 411226 3732
rect 428458 3720 428464 3732
rect 411220 3692 428464 3720
rect 411220 3680 411226 3692
rect 428458 3680 428464 3692
rect 428516 3680 428522 3732
rect 431770 3680 431776 3732
rect 431828 3720 431834 3732
rect 450906 3720 450912 3732
rect 431828 3692 450912 3720
rect 431828 3680 431834 3692
rect 450906 3680 450912 3692
rect 450964 3680 450970 3732
rect 452470 3680 452476 3732
rect 452528 3720 452534 3732
rect 453761 3723 453819 3729
rect 453761 3720 453773 3723
rect 452528 3692 453773 3720
rect 452528 3680 452534 3692
rect 453761 3689 453773 3692
rect 453807 3689 453819 3723
rect 453761 3683 453819 3689
rect 453942 3680 453948 3732
rect 454000 3720 454006 3732
rect 474550 3720 474556 3732
rect 454000 3692 474556 3720
rect 454000 3680 454006 3692
rect 474550 3680 474556 3692
rect 474608 3680 474614 3732
rect 474642 3680 474648 3732
rect 474700 3720 474706 3732
rect 495894 3720 495900 3732
rect 474700 3692 495900 3720
rect 474700 3680 474706 3692
rect 495894 3680 495900 3692
rect 495952 3680 495958 3732
rect 496722 3680 496728 3732
rect 496780 3720 496786 3732
rect 520734 3720 520740 3732
rect 496780 3692 520740 3720
rect 496780 3680 496786 3692
rect 520734 3680 520740 3692
rect 520792 3680 520798 3732
rect 526990 3680 526996 3732
rect 527048 3720 527054 3732
rect 552658 3720 552664 3732
rect 527048 3692 552664 3720
rect 527048 3680 527054 3692
rect 552658 3680 552664 3692
rect 552716 3680 552722 3732
rect 553302 3680 553308 3732
rect 553360 3720 553366 3732
rect 582190 3720 582196 3732
rect 553360 3692 582196 3720
rect 553360 3680 553366 3692
rect 582190 3680 582196 3692
rect 582248 3680 582254 3732
rect 371694 3652 371700 3664
rect 358832 3624 371700 3652
rect 371694 3612 371700 3624
rect 371752 3612 371758 3664
rect 375282 3612 375288 3664
rect 375340 3652 375346 3664
rect 389450 3652 389456 3664
rect 375340 3624 389456 3652
rect 375340 3612 375346 3624
rect 389450 3612 389456 3624
rect 389508 3612 389514 3664
rect 390462 3612 390468 3664
rect 390520 3652 390526 3664
rect 406010 3652 406016 3664
rect 390520 3624 406016 3652
rect 390520 3612 390526 3624
rect 406010 3612 406016 3624
rect 406068 3612 406074 3664
rect 407022 3612 407028 3664
rect 407080 3652 407086 3664
rect 423766 3652 423772 3664
rect 407080 3624 423772 3652
rect 407080 3612 407086 3624
rect 423766 3612 423772 3624
rect 423824 3612 423830 3664
rect 427722 3612 427728 3664
rect 427780 3652 427786 3664
rect 446214 3652 446220 3664
rect 427780 3624 446220 3652
rect 427780 3612 427786 3624
rect 446214 3612 446220 3624
rect 446272 3612 446278 3664
rect 448330 3612 448336 3664
rect 448388 3652 448394 3664
rect 468662 3652 468668 3664
rect 448388 3624 468668 3652
rect 448388 3612 448394 3624
rect 468662 3612 468668 3624
rect 468720 3612 468726 3664
rect 474458 3612 474464 3664
rect 474516 3652 474522 3664
rect 497090 3652 497096 3664
rect 474516 3624 497096 3652
rect 474516 3612 474522 3624
rect 497090 3612 497096 3624
rect 497148 3612 497154 3664
rect 498102 3612 498108 3664
rect 498160 3652 498166 3664
rect 521838 3652 521844 3664
rect 498160 3624 521844 3652
rect 498160 3612 498166 3624
rect 521838 3612 521844 3624
rect 521896 3612 521902 3664
rect 522942 3612 522948 3664
rect 523000 3652 523006 3664
rect 549070 3652 549076 3664
rect 523000 3624 549076 3652
rect 523000 3612 523006 3624
rect 549070 3612 549076 3624
rect 549128 3612 549134 3664
rect 550542 3612 550548 3664
rect 550600 3652 550606 3664
rect 578602 3652 578608 3664
rect 550600 3624 578608 3652
rect 550600 3612 550606 3624
rect 578602 3612 578608 3624
rect 578660 3612 578666 3664
rect 338022 3544 338028 3596
rect 338080 3584 338086 3596
rect 349246 3584 349252 3596
rect 338080 3556 349252 3584
rect 338080 3544 338086 3556
rect 349246 3544 349252 3556
rect 349304 3544 349310 3596
rect 353202 3544 353208 3596
rect 353260 3584 353266 3596
rect 365806 3584 365812 3596
rect 353260 3556 365812 3584
rect 353260 3544 353266 3556
rect 365806 3544 365812 3556
rect 365864 3544 365870 3596
rect 368290 3544 368296 3596
rect 368348 3584 368354 3596
rect 381170 3584 381176 3596
rect 368348 3556 381176 3584
rect 368348 3544 368354 3556
rect 381170 3544 381176 3556
rect 381228 3544 381234 3596
rect 383562 3544 383568 3596
rect 383620 3584 383626 3596
rect 398926 3584 398932 3596
rect 383620 3556 398932 3584
rect 383620 3544 383626 3556
rect 398926 3544 398932 3556
rect 398984 3544 398990 3596
rect 400030 3544 400036 3596
rect 400088 3584 400094 3596
rect 415486 3584 415492 3596
rect 400088 3556 415492 3584
rect 400088 3544 400094 3556
rect 415486 3544 415492 3556
rect 415544 3544 415550 3596
rect 420822 3544 420828 3596
rect 420880 3584 420886 3596
rect 439130 3584 439136 3596
rect 420880 3556 439136 3584
rect 420880 3544 420886 3556
rect 439130 3544 439136 3556
rect 439188 3544 439194 3596
rect 442810 3544 442816 3596
rect 442868 3584 442874 3596
rect 462774 3584 462780 3596
rect 442868 3556 462780 3584
rect 442868 3544 442874 3556
rect 462774 3544 462780 3556
rect 462832 3544 462838 3596
rect 464982 3544 464988 3596
rect 465040 3584 465046 3596
rect 486418 3584 486424 3596
rect 465040 3556 486424 3584
rect 465040 3544 465046 3556
rect 486418 3544 486424 3556
rect 486476 3544 486482 3596
rect 489822 3544 489828 3596
rect 489880 3584 489886 3596
rect 513558 3584 513564 3596
rect 489880 3556 513564 3584
rect 489880 3544 489886 3556
rect 513558 3544 513564 3556
rect 513616 3544 513622 3596
rect 520182 3544 520188 3596
rect 520240 3584 520246 3596
rect 545482 3584 545488 3596
rect 520240 3556 545488 3584
rect 520240 3544 520246 3556
rect 545482 3544 545488 3556
rect 545540 3544 545546 3596
rect 549162 3544 549168 3596
rect 549220 3584 549226 3596
rect 577406 3584 577412 3596
rect 549220 3556 577412 3584
rect 549220 3544 549226 3556
rect 577406 3544 577412 3556
rect 577464 3544 577470 3596
rect 342162 3516 342168 3528
rect 332796 3488 342168 3516
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 344922 3476 344928 3528
rect 344980 3516 344986 3528
rect 356330 3516 356336 3528
rect 344980 3488 356336 3516
rect 344980 3476 344986 3488
rect 356330 3476 356336 3488
rect 356388 3476 356394 3528
rect 358633 3519 358691 3525
rect 358633 3485 358645 3519
rect 358679 3516 358691 3519
rect 361114 3516 361120 3528
rect 358679 3488 361120 3516
rect 358679 3485 358691 3488
rect 358633 3479 358691 3485
rect 361114 3476 361120 3488
rect 361172 3476 361178 3528
rect 370590 3516 370596 3528
rect 361316 3488 370596 3516
rect 73798 3408 73804 3460
rect 73856 3448 73862 3460
rect 74442 3448 74448 3460
rect 73856 3420 74448 3448
rect 73856 3408 73862 3420
rect 74442 3408 74448 3420
rect 74500 3408 74506 3460
rect 131758 3408 131764 3460
rect 131816 3448 131822 3460
rect 132402 3448 132408 3460
rect 131816 3420 132408 3448
rect 131816 3408 131822 3420
rect 132402 3408 132408 3420
rect 132460 3408 132466 3460
rect 135254 3408 135260 3460
rect 135312 3448 135318 3460
rect 136542 3448 136548 3460
rect 135312 3420 136548 3448
rect 135312 3408 135318 3420
rect 136542 3408 136548 3420
rect 136600 3408 136606 3460
rect 155402 3408 155408 3460
rect 155460 3448 155466 3460
rect 155862 3448 155868 3460
rect 155460 3420 155868 3448
rect 155460 3408 155466 3420
rect 155862 3408 155868 3420
rect 155920 3408 155926 3460
rect 195974 3408 195980 3460
rect 196032 3448 196038 3460
rect 196802 3448 196808 3460
rect 196032 3420 196808 3448
rect 196032 3408 196038 3420
rect 196802 3408 196808 3420
rect 196860 3408 196866 3460
rect 216582 3408 216588 3460
rect 216640 3448 216646 3460
rect 218054 3448 218060 3460
rect 216640 3420 218060 3448
rect 216640 3408 216646 3420
rect 218054 3408 218060 3420
rect 218112 3408 218118 3460
rect 224862 3408 224868 3460
rect 224920 3448 224926 3460
rect 227530 3448 227536 3460
rect 224920 3420 227536 3448
rect 224920 3408 224926 3420
rect 227530 3408 227536 3420
rect 227588 3408 227594 3460
rect 231762 3408 231768 3460
rect 231820 3448 231826 3460
rect 234614 3448 234620 3460
rect 231820 3420 234620 3448
rect 231820 3408 231826 3420
rect 234614 3408 234620 3420
rect 234672 3408 234678 3460
rect 241422 3408 241428 3460
rect 241480 3448 241486 3460
rect 245194 3448 245200 3460
rect 241480 3420 245200 3448
rect 241480 3408 241486 3420
rect 245194 3408 245200 3420
rect 245252 3408 245258 3460
rect 249702 3408 249708 3460
rect 249760 3448 249766 3460
rect 253474 3448 253480 3460
rect 249760 3420 253480 3448
rect 249760 3408 249766 3420
rect 253474 3408 253480 3420
rect 253532 3408 253538 3460
rect 259362 3408 259368 3460
rect 259420 3448 259426 3460
rect 264146 3448 264152 3460
rect 259420 3420 264152 3448
rect 259420 3408 259426 3420
rect 264146 3408 264152 3420
rect 264204 3408 264210 3460
rect 267550 3408 267556 3460
rect 267608 3448 267614 3460
rect 273622 3448 273628 3460
rect 267608 3420 273628 3448
rect 267608 3408 267614 3420
rect 273622 3408 273628 3420
rect 273680 3408 273686 3460
rect 277210 3408 277216 3460
rect 277268 3448 277274 3460
rect 284294 3448 284300 3460
rect 277268 3420 284300 3448
rect 277268 3408 277274 3420
rect 284294 3408 284300 3420
rect 284352 3408 284358 3460
rect 296622 3408 296628 3460
rect 296680 3448 296686 3460
rect 304350 3448 304356 3460
rect 296680 3420 304356 3448
rect 296680 3408 296686 3420
rect 304350 3408 304356 3420
rect 304408 3408 304414 3460
rect 304810 3408 304816 3460
rect 304868 3448 304874 3460
rect 313826 3448 313832 3460
rect 304868 3420 313832 3448
rect 304868 3408 304874 3420
rect 313826 3408 313832 3420
rect 313884 3408 313890 3460
rect 314470 3408 314476 3460
rect 314528 3448 314534 3460
rect 324406 3448 324412 3460
rect 314528 3420 324412 3448
rect 314528 3408 314534 3420
rect 324406 3408 324412 3420
rect 324464 3408 324470 3460
rect 325694 3408 325700 3460
rect 325752 3448 325758 3460
rect 336274 3448 336280 3460
rect 325752 3420 336280 3448
rect 325752 3408 325758 3420
rect 336274 3408 336280 3420
rect 336332 3408 336338 3460
rect 336550 3408 336556 3460
rect 336608 3448 336614 3460
rect 348050 3448 348056 3460
rect 336608 3420 348056 3448
rect 336608 3408 336614 3420
rect 348050 3408 348056 3420
rect 348108 3408 348114 3460
rect 351822 3408 351828 3460
rect 351880 3448 351886 3460
rect 361209 3451 361267 3457
rect 361209 3448 361221 3451
rect 351880 3420 361221 3448
rect 351880 3408 351886 3420
rect 361209 3417 361221 3420
rect 361255 3417 361267 3451
rect 361209 3411 361267 3417
rect 300670 3340 300676 3392
rect 300728 3380 300734 3392
rect 309042 3380 309048 3392
rect 300728 3352 309048 3380
rect 300728 3340 300734 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 319990 3340 319996 3392
rect 320048 3380 320054 3392
rect 330386 3380 330392 3392
rect 320048 3352 330392 3380
rect 320048 3340 320054 3352
rect 330386 3340 330392 3352
rect 330444 3340 330450 3392
rect 333790 3340 333796 3392
rect 333848 3380 333854 3392
rect 344554 3380 344560 3392
rect 333848 3352 344560 3380
rect 333848 3340 333854 3352
rect 344554 3340 344560 3352
rect 344612 3340 344618 3392
rect 357250 3340 357256 3392
rect 357308 3380 357314 3392
rect 361316 3380 361344 3488
rect 370590 3476 370596 3488
rect 370648 3476 370654 3528
rect 379330 3476 379336 3528
rect 379388 3516 379394 3528
rect 394234 3516 394240 3528
rect 379388 3488 394240 3516
rect 379388 3476 379394 3488
rect 394234 3476 394240 3488
rect 394292 3476 394298 3528
rect 397362 3476 397368 3528
rect 397420 3516 397426 3528
rect 413094 3516 413100 3528
rect 397420 3488 413100 3516
rect 397420 3476 397426 3488
rect 413094 3476 413100 3488
rect 413152 3476 413158 3528
rect 415210 3476 415216 3528
rect 415268 3516 415274 3528
rect 433242 3516 433248 3528
rect 415268 3488 433248 3516
rect 415268 3476 415274 3488
rect 433242 3476 433248 3488
rect 433300 3476 433306 3528
rect 437382 3476 437388 3528
rect 437440 3516 437446 3528
rect 456886 3516 456892 3528
rect 437440 3488 456892 3516
rect 437440 3476 437446 3488
rect 456886 3476 456892 3488
rect 456944 3476 456950 3528
rect 458082 3476 458088 3528
rect 458140 3516 458146 3528
rect 479334 3516 479340 3528
rect 458140 3488 479340 3516
rect 458140 3476 458146 3488
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 480162 3476 480168 3528
rect 480220 3516 480226 3528
rect 502978 3516 502984 3528
rect 480220 3488 502984 3516
rect 480220 3476 480226 3488
rect 502978 3476 502984 3488
rect 503036 3476 503042 3528
rect 506382 3476 506388 3528
rect 506440 3516 506446 3528
rect 531314 3516 531320 3528
rect 506440 3488 531320 3516
rect 506440 3476 506446 3488
rect 531314 3476 531320 3488
rect 531372 3476 531378 3528
rect 543550 3476 543556 3528
rect 543608 3516 543614 3528
rect 571518 3516 571524 3528
rect 543608 3488 571524 3516
rect 543608 3476 543614 3488
rect 571518 3476 571524 3488
rect 571576 3476 571582 3528
rect 361393 3451 361451 3457
rect 361393 3417 361405 3451
rect 361439 3448 361451 3451
rect 364610 3448 364616 3460
rect 361439 3420 364616 3448
rect 361439 3417 361451 3420
rect 361393 3411 361451 3417
rect 364610 3408 364616 3420
rect 364668 3408 364674 3460
rect 368382 3408 368388 3460
rect 368440 3448 368446 3460
rect 382366 3448 382372 3460
rect 368440 3420 382372 3448
rect 368440 3408 368446 3420
rect 382366 3408 382372 3420
rect 382424 3408 382430 3460
rect 388990 3408 388996 3460
rect 389048 3448 389054 3460
rect 404814 3448 404820 3460
rect 389048 3420 404820 3448
rect 389048 3408 389054 3420
rect 404814 3408 404820 3420
rect 404872 3408 404878 3460
rect 405550 3408 405556 3460
rect 405608 3448 405614 3460
rect 422570 3448 422576 3460
rect 405608 3420 422576 3448
rect 405608 3408 405614 3420
rect 422570 3408 422576 3420
rect 422628 3408 422634 3460
rect 426250 3408 426256 3460
rect 426308 3448 426314 3460
rect 445018 3448 445024 3460
rect 426308 3420 445024 3448
rect 426308 3408 426314 3420
rect 445018 3408 445024 3420
rect 445076 3408 445082 3460
rect 449894 3408 449900 3460
rect 449952 3448 449958 3460
rect 453761 3451 453819 3457
rect 449952 3420 453712 3448
rect 449952 3408 449958 3420
rect 369394 3380 369400 3392
rect 357308 3352 361344 3380
rect 362420 3352 369400 3380
rect 357308 3340 357314 3352
rect 80882 3272 80888 3324
rect 80940 3312 80946 3324
rect 81342 3312 81348 3324
rect 80940 3284 81348 3312
rect 80940 3272 80946 3284
rect 81342 3272 81348 3284
rect 81400 3272 81406 3324
rect 85666 3272 85672 3324
rect 85724 3312 85730 3324
rect 86770 3312 86776 3324
rect 85724 3284 86776 3312
rect 85724 3272 85730 3284
rect 86770 3272 86776 3284
rect 86828 3272 86834 3324
rect 89162 3272 89168 3324
rect 89220 3312 89226 3324
rect 89622 3312 89628 3324
rect 89220 3284 89628 3312
rect 89220 3272 89226 3284
rect 89622 3272 89628 3284
rect 89680 3272 89686 3324
rect 126974 3272 126980 3324
rect 127032 3312 127038 3324
rect 130378 3312 130384 3324
rect 127032 3284 130384 3312
rect 127032 3272 127038 3284
rect 130378 3272 130384 3284
rect 130436 3272 130442 3324
rect 220722 3272 220728 3324
rect 220780 3312 220786 3324
rect 222746 3312 222752 3324
rect 220780 3284 222752 3312
rect 220780 3272 220786 3284
rect 222746 3272 222752 3284
rect 222804 3272 222810 3324
rect 252462 3272 252468 3324
rect 252520 3312 252526 3324
rect 257062 3312 257068 3324
rect 252520 3284 257068 3312
rect 252520 3272 252526 3284
rect 257062 3272 257068 3284
rect 257120 3272 257126 3324
rect 260742 3272 260748 3324
rect 260800 3312 260806 3324
rect 265342 3312 265348 3324
rect 260800 3284 265348 3312
rect 260800 3272 260806 3284
rect 265342 3272 265348 3284
rect 265400 3272 265406 3324
rect 271782 3272 271788 3324
rect 271840 3312 271846 3324
rect 277118 3312 277124 3324
rect 271840 3284 277124 3312
rect 271840 3272 271846 3284
rect 277118 3272 277124 3284
rect 277176 3272 277182 3324
rect 278682 3272 278688 3324
rect 278740 3312 278746 3324
rect 285398 3312 285404 3324
rect 278740 3284 285404 3312
rect 278740 3272 278746 3284
rect 285398 3272 285404 3284
rect 285456 3272 285462 3324
rect 288250 3272 288256 3324
rect 288308 3312 288314 3324
rect 296070 3312 296076 3324
rect 288308 3284 296076 3312
rect 288308 3272 288314 3284
rect 296070 3272 296076 3284
rect 296128 3272 296134 3324
rect 298002 3272 298008 3324
rect 298060 3312 298066 3324
rect 305546 3312 305552 3324
rect 298060 3284 305552 3312
rect 298060 3272 298066 3284
rect 305546 3272 305552 3284
rect 305604 3272 305610 3324
rect 350350 3272 350356 3324
rect 350408 3312 350414 3324
rect 362310 3312 362316 3324
rect 350408 3284 362316 3312
rect 350408 3272 350414 3284
rect 362310 3272 362316 3284
rect 362368 3272 362374 3324
rect 84470 3204 84476 3256
rect 84528 3244 84534 3256
rect 85482 3244 85488 3256
rect 84528 3216 85488 3244
rect 84528 3204 84534 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 208302 3204 208308 3256
rect 208360 3244 208366 3256
rect 209774 3244 209780 3256
rect 208360 3216 209780 3244
rect 208360 3204 208366 3216
rect 209774 3204 209780 3216
rect 209832 3204 209838 3256
rect 245562 3204 245568 3256
rect 245620 3244 245626 3256
rect 245620 3216 248414 3244
rect 245620 3204 245626 3216
rect 230382 3136 230388 3188
rect 230440 3176 230446 3188
rect 233418 3176 233424 3188
rect 230440 3148 233424 3176
rect 230440 3136 230446 3148
rect 233418 3136 233424 3148
rect 233476 3136 233482 3188
rect 234522 3136 234528 3188
rect 234580 3176 234586 3188
rect 237006 3176 237012 3188
rect 234580 3148 237012 3176
rect 234580 3136 234586 3148
rect 237006 3136 237012 3148
rect 237064 3136 237070 3188
rect 240042 3136 240048 3188
rect 240100 3176 240106 3188
rect 242894 3176 242900 3188
rect 240100 3148 242900 3176
rect 240100 3136 240106 3148
rect 242894 3136 242900 3148
rect 242952 3136 242958 3188
rect 246298 3136 246304 3188
rect 246356 3176 246362 3188
rect 247586 3176 247592 3188
rect 246356 3148 247592 3176
rect 246356 3136 246362 3148
rect 247586 3136 247592 3148
rect 247644 3136 247650 3188
rect 248386 3176 248414 3216
rect 250990 3204 250996 3256
rect 251048 3244 251054 3256
rect 254670 3244 254676 3256
rect 251048 3216 254676 3244
rect 251048 3204 251054 3216
rect 254670 3204 254676 3216
rect 254728 3204 254734 3256
rect 340782 3204 340788 3256
rect 340840 3244 340846 3256
rect 351638 3244 351644 3256
rect 340840 3216 351644 3244
rect 340840 3204 340846 3216
rect 351638 3204 351644 3216
rect 351696 3204 351702 3256
rect 357342 3204 357348 3256
rect 357400 3244 357406 3256
rect 362420 3244 362448 3352
rect 369394 3340 369400 3352
rect 369452 3340 369458 3392
rect 372522 3340 372528 3392
rect 372580 3380 372586 3392
rect 385954 3380 385960 3392
rect 372580 3352 385960 3380
rect 372580 3340 372586 3352
rect 385954 3340 385960 3352
rect 386012 3340 386018 3392
rect 386322 3340 386328 3392
rect 386380 3380 386386 3392
rect 401318 3380 401324 3392
rect 386380 3352 401324 3380
rect 386380 3340 386386 3352
rect 401318 3340 401324 3352
rect 401376 3340 401382 3392
rect 405568 3352 408816 3380
rect 364242 3272 364248 3324
rect 364300 3312 364306 3324
rect 377674 3312 377680 3324
rect 364300 3284 377680 3312
rect 364300 3272 364306 3284
rect 377674 3272 377680 3284
rect 377732 3272 377738 3324
rect 389082 3272 389088 3324
rect 389140 3312 389146 3324
rect 403618 3312 403624 3324
rect 389140 3284 403624 3312
rect 389140 3272 389146 3284
rect 403618 3272 403624 3284
rect 403676 3272 403682 3324
rect 357400 3216 362448 3244
rect 357400 3204 357406 3216
rect 362862 3204 362868 3256
rect 362920 3244 362926 3256
rect 375282 3244 375288 3256
rect 362920 3216 375288 3244
rect 362920 3204 362926 3216
rect 375282 3204 375288 3216
rect 375340 3204 375346 3256
rect 379422 3204 379428 3256
rect 379480 3244 379486 3256
rect 393038 3244 393044 3256
rect 379480 3216 393044 3244
rect 379480 3204 379486 3216
rect 393038 3204 393044 3216
rect 393096 3204 393102 3256
rect 401502 3204 401508 3256
rect 401560 3244 401566 3256
rect 405568 3244 405596 3352
rect 405642 3272 405648 3324
rect 405700 3312 405706 3324
rect 405700 3284 408724 3312
rect 405700 3272 405706 3284
rect 401560 3216 405596 3244
rect 401560 3204 401566 3216
rect 248782 3176 248788 3188
rect 248386 3148 248788 3176
rect 248782 3136 248788 3148
rect 248840 3136 248846 3188
rect 264238 3136 264244 3188
rect 264296 3176 264302 3188
rect 266538 3176 266544 3188
rect 264296 3148 266544 3176
rect 264296 3136 264302 3148
rect 266538 3136 266544 3148
rect 266596 3136 266602 3188
rect 273162 3136 273168 3188
rect 273220 3176 273226 3188
rect 279510 3176 279516 3188
rect 273220 3148 279516 3176
rect 273220 3136 273226 3148
rect 279510 3136 279516 3148
rect 279568 3136 279574 3188
rect 369762 3136 369768 3188
rect 369820 3176 369826 3188
rect 383562 3176 383568 3188
rect 369820 3148 383568 3176
rect 369820 3136 369826 3148
rect 383562 3136 383568 3148
rect 383620 3136 383626 3188
rect 387702 3136 387708 3188
rect 387760 3176 387766 3188
rect 402514 3176 402520 3188
rect 387760 3148 402520 3176
rect 387760 3136 387766 3148
rect 402514 3136 402520 3148
rect 402572 3136 402578 3188
rect 408310 3136 408316 3188
rect 408368 3176 408374 3188
rect 408696 3176 408724 3284
rect 408788 3244 408816 3352
rect 413922 3340 413928 3392
rect 413980 3380 413986 3392
rect 430850 3380 430856 3392
rect 413980 3352 430856 3380
rect 413980 3340 413986 3352
rect 430850 3340 430856 3352
rect 430908 3340 430914 3392
rect 445662 3340 445668 3392
rect 445720 3380 445726 3392
rect 445720 3352 449848 3380
rect 445720 3340 445726 3352
rect 409782 3272 409788 3324
rect 409840 3312 409846 3324
rect 426158 3312 426164 3324
rect 409840 3284 426164 3312
rect 409840 3272 409846 3284
rect 426158 3272 426164 3284
rect 426216 3272 426222 3324
rect 431862 3272 431868 3324
rect 431920 3312 431926 3324
rect 449710 3312 449716 3324
rect 431920 3284 449716 3312
rect 431920 3272 431926 3284
rect 449710 3272 449716 3284
rect 449768 3272 449774 3324
rect 449820 3312 449848 3352
rect 453577 3315 453635 3321
rect 453577 3312 453589 3315
rect 449820 3284 453589 3312
rect 453577 3281 453589 3284
rect 453623 3281 453635 3315
rect 453684 3312 453712 3420
rect 453761 3417 453773 3451
rect 453807 3448 453819 3451
rect 473446 3448 473452 3460
rect 453807 3420 473452 3448
rect 453807 3417 453819 3420
rect 453761 3411 453819 3417
rect 473446 3408 473452 3420
rect 473504 3408 473510 3460
rect 491202 3408 491208 3460
rect 491260 3448 491266 3460
rect 514754 3448 514760 3460
rect 491260 3420 514760 3448
rect 491260 3408 491266 3420
rect 514754 3408 514760 3420
rect 514812 3408 514818 3460
rect 517330 3408 517336 3460
rect 517388 3448 517394 3460
rect 543182 3448 543188 3460
rect 517388 3420 543188 3448
rect 517388 3408 517394 3420
rect 543182 3408 543188 3420
rect 543240 3408 543246 3460
rect 551922 3408 551928 3460
rect 551980 3448 551986 3460
rect 580994 3448 581000 3460
rect 551980 3420 581000 3448
rect 551980 3408 551986 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 453853 3383 453911 3389
rect 453853 3349 453865 3383
rect 453899 3380 453911 3383
rect 465166 3380 465172 3392
rect 453899 3352 465172 3380
rect 453899 3349 453911 3352
rect 453853 3343 453911 3349
rect 465166 3340 465172 3352
rect 465224 3340 465230 3392
rect 469122 3340 469128 3392
rect 469180 3380 469186 3392
rect 489914 3380 489920 3392
rect 469180 3352 489920 3380
rect 469180 3340 469186 3352
rect 489914 3340 489920 3352
rect 489972 3340 489978 3392
rect 500862 3340 500868 3392
rect 500920 3380 500926 3392
rect 525426 3380 525432 3392
rect 500920 3352 525432 3380
rect 500920 3340 500926 3352
rect 525426 3340 525432 3352
rect 525484 3340 525490 3392
rect 527082 3340 527088 3392
rect 527140 3380 527146 3392
rect 553762 3380 553768 3392
rect 527140 3352 553768 3380
rect 527140 3340 527146 3352
rect 553762 3340 553768 3352
rect 553820 3340 553826 3392
rect 469858 3312 469864 3324
rect 453684 3284 469864 3312
rect 453577 3275 453635 3281
rect 469858 3272 469864 3284
rect 469916 3272 469922 3324
rect 471882 3272 471888 3324
rect 471940 3312 471946 3324
rect 493502 3312 493508 3324
rect 471940 3284 493508 3312
rect 471940 3272 471946 3284
rect 493502 3272 493508 3284
rect 493560 3272 493566 3324
rect 503622 3272 503628 3324
rect 503680 3312 503686 3324
rect 527818 3312 527824 3324
rect 503680 3284 527824 3312
rect 503680 3272 503686 3284
rect 527818 3272 527824 3284
rect 527876 3272 527882 3324
rect 532602 3272 532608 3324
rect 532660 3312 532666 3324
rect 559742 3312 559748 3324
rect 532660 3284 559748 3312
rect 532660 3272 532666 3284
rect 559742 3272 559748 3284
rect 559800 3272 559806 3324
rect 417878 3244 417884 3256
rect 408788 3216 417884 3244
rect 417878 3204 417884 3216
rect 417936 3204 417942 3256
rect 418062 3204 418068 3256
rect 418120 3244 418126 3256
rect 435542 3244 435548 3256
rect 418120 3216 435548 3244
rect 418120 3204 418126 3216
rect 435542 3204 435548 3216
rect 435600 3204 435606 3256
rect 440142 3204 440148 3256
rect 440200 3244 440206 3256
rect 459186 3244 459192 3256
rect 440200 3216 459192 3244
rect 440200 3204 440206 3216
rect 459186 3204 459192 3216
rect 459244 3204 459250 3256
rect 462222 3204 462228 3256
rect 462280 3244 462286 3256
rect 482830 3244 482836 3256
rect 462280 3216 482836 3244
rect 462280 3204 462286 3216
rect 482830 3204 482836 3216
rect 482888 3204 482894 3256
rect 488442 3204 488448 3256
rect 488500 3244 488506 3256
rect 511258 3244 511264 3256
rect 488500 3216 511264 3244
rect 488500 3204 488506 3216
rect 511258 3204 511264 3216
rect 511316 3204 511322 3256
rect 511902 3204 511908 3256
rect 511960 3244 511966 3256
rect 536098 3244 536104 3256
rect 511960 3216 536104 3244
rect 511960 3204 511966 3216
rect 536098 3204 536104 3216
rect 536156 3204 536162 3256
rect 536742 3204 536748 3256
rect 536800 3244 536806 3256
rect 563238 3244 563244 3256
rect 536800 3216 563244 3244
rect 536800 3204 536806 3216
rect 563238 3204 563244 3216
rect 563296 3204 563302 3256
rect 421374 3176 421380 3188
rect 408368 3148 408540 3176
rect 408696 3148 421380 3176
rect 408368 3136 408374 3148
rect 378042 3068 378048 3120
rect 378100 3108 378106 3120
rect 391842 3108 391848 3120
rect 378100 3080 391848 3108
rect 378100 3068 378106 3080
rect 391842 3068 391848 3080
rect 391900 3068 391906 3120
rect 393222 3068 393228 3120
rect 393280 3108 393286 3120
rect 408402 3108 408408 3120
rect 393280 3080 408408 3108
rect 393280 3068 393286 3080
rect 408402 3068 408408 3080
rect 408460 3068 408466 3120
rect 408512 3108 408540 3148
rect 421374 3136 421380 3148
rect 421432 3136 421438 3188
rect 424870 3136 424876 3188
rect 424928 3176 424934 3188
rect 424928 3148 431954 3176
rect 424928 3136 424934 3148
rect 424962 3108 424968 3120
rect 408512 3080 424968 3108
rect 424962 3068 424968 3080
rect 425020 3068 425026 3120
rect 431926 3108 431954 3148
rect 433150 3136 433156 3188
rect 433208 3176 433214 3188
rect 452102 3176 452108 3188
rect 433208 3148 452108 3176
rect 433208 3136 433214 3148
rect 452102 3136 452108 3148
rect 452160 3136 452166 3188
rect 452562 3136 452568 3188
rect 452620 3176 452626 3188
rect 454589 3179 454647 3185
rect 454589 3176 454601 3179
rect 452620 3148 454601 3176
rect 452620 3136 452626 3148
rect 454589 3145 454601 3148
rect 454635 3145 454647 3179
rect 454589 3139 454647 3145
rect 455322 3136 455328 3188
rect 455380 3176 455386 3188
rect 475746 3176 475752 3188
rect 455380 3148 475752 3176
rect 455380 3136 455386 3148
rect 475746 3136 475752 3148
rect 475804 3136 475810 3188
rect 478782 3136 478788 3188
rect 478840 3176 478846 3188
rect 500586 3176 500592 3188
rect 478840 3148 500592 3176
rect 478840 3136 478846 3148
rect 500586 3136 500592 3148
rect 500644 3136 500650 3188
rect 517422 3136 517428 3188
rect 517480 3176 517486 3188
rect 541986 3176 541992 3188
rect 517480 3148 541992 3176
rect 517480 3136 517486 3148
rect 541986 3136 541992 3148
rect 542044 3136 542050 3188
rect 547782 3136 547788 3188
rect 547840 3176 547846 3188
rect 575106 3176 575112 3188
rect 547840 3148 575112 3176
rect 547840 3136 547846 3148
rect 575106 3136 575112 3148
rect 575164 3136 575170 3188
rect 442626 3108 442632 3120
rect 431926 3080 442632 3108
rect 442626 3068 442632 3080
rect 442684 3068 442690 3120
rect 448422 3068 448428 3120
rect 448480 3108 448486 3120
rect 467466 3108 467472 3120
rect 448480 3080 467472 3108
rect 448480 3068 448486 3080
rect 467466 3068 467472 3080
rect 467524 3068 467530 3120
rect 467742 3068 467748 3120
rect 467800 3108 467806 3120
rect 488810 3108 488816 3120
rect 467800 3080 488816 3108
rect 467800 3068 467806 3080
rect 488810 3068 488816 3080
rect 488868 3068 488874 3120
rect 500770 3068 500776 3120
rect 500828 3108 500834 3120
rect 524230 3108 524236 3120
rect 500828 3080 524236 3108
rect 500828 3068 500834 3080
rect 524230 3068 524236 3080
rect 524288 3068 524294 3120
rect 540882 3068 540888 3120
rect 540940 3108 540946 3120
rect 568022 3108 568028 3120
rect 540940 3080 568028 3108
rect 540940 3068 540946 3080
rect 568022 3068 568028 3080
rect 568080 3068 568086 3120
rect 143534 3000 143540 3052
rect 143592 3040 143598 3052
rect 144638 3040 144644 3052
rect 143592 3012 144644 3040
rect 143592 3000 143598 3012
rect 144638 3000 144644 3012
rect 144696 3000 144702 3052
rect 150618 3000 150624 3052
rect 150676 3040 150682 3052
rect 151722 3040 151728 3052
rect 150676 3012 151728 3040
rect 150676 3000 150682 3012
rect 151722 3000 151728 3012
rect 151780 3000 151786 3052
rect 263502 3000 263508 3052
rect 263560 3040 263566 3052
rect 268838 3040 268844 3052
rect 263560 3012 268844 3040
rect 263560 3000 263566 3012
rect 268838 3000 268844 3012
rect 268896 3000 268902 3052
rect 291102 3000 291108 3052
rect 291160 3040 291166 3052
rect 298462 3040 298468 3052
rect 291160 3012 298468 3040
rect 291160 3000 291166 3012
rect 298462 3000 298468 3012
rect 298520 3000 298526 3052
rect 402882 3000 402888 3052
rect 402940 3040 402946 3052
rect 418982 3040 418988 3052
rect 402940 3012 418988 3040
rect 402940 3000 402946 3012
rect 418982 3000 418988 3012
rect 419040 3000 419046 3052
rect 419442 3000 419448 3052
rect 419500 3040 419506 3052
rect 436738 3040 436744 3052
rect 419500 3012 436744 3040
rect 419500 3000 419506 3012
rect 436738 3000 436744 3012
rect 436796 3000 436802 3052
rect 438762 3000 438768 3052
rect 438820 3040 438826 3052
rect 458082 3040 458088 3052
rect 438820 3012 458088 3040
rect 438820 3000 438826 3012
rect 458082 3000 458088 3012
rect 458140 3000 458146 3052
rect 495342 3000 495348 3052
rect 495400 3040 495406 3052
rect 518342 3040 518348 3052
rect 495400 3012 518348 3040
rect 495400 3000 495406 3012
rect 518342 3000 518348 3012
rect 518400 3000 518406 3052
rect 538122 3000 538128 3052
rect 538180 3040 538186 3052
rect 564434 3040 564440 3052
rect 538180 3012 564440 3040
rect 538180 3000 538186 3012
rect 564434 3000 564440 3012
rect 564492 3000 564498 3052
rect 582377 3043 582435 3049
rect 582377 3009 582389 3043
rect 582423 3040 582435 3043
rect 583386 3040 583392 3052
rect 582423 3012 583392 3040
rect 582423 3009 582435 3012
rect 582377 3003 582435 3009
rect 583386 3000 583392 3012
rect 583444 3000 583450 3052
rect 25314 2932 25320 2984
rect 25372 2972 25378 2984
rect 26142 2972 26148 2984
rect 25372 2944 26148 2972
rect 25372 2932 25378 2944
rect 26142 2932 26148 2944
rect 26200 2932 26206 2984
rect 83274 2932 83280 2984
rect 83332 2972 83338 2984
rect 84102 2972 84108 2984
rect 83332 2944 84108 2972
rect 83332 2932 83338 2944
rect 84102 2932 84108 2944
rect 84160 2932 84166 2984
rect 213822 2932 213828 2984
rect 213880 2972 213886 2984
rect 215662 2972 215668 2984
rect 213880 2944 215668 2972
rect 213880 2932 213886 2944
rect 215662 2932 215668 2944
rect 215720 2932 215726 2984
rect 224770 2932 224776 2984
rect 224828 2972 224834 2984
rect 226334 2972 226340 2984
rect 224828 2944 226340 2972
rect 224828 2932 224834 2944
rect 226334 2932 226340 2944
rect 226392 2932 226398 2984
rect 270402 2932 270408 2984
rect 270460 2972 270466 2984
rect 276014 2972 276020 2984
rect 270460 2944 276020 2972
rect 270460 2932 270466 2944
rect 276014 2932 276020 2944
rect 276072 2932 276078 2984
rect 280062 2932 280068 2984
rect 280120 2972 280126 2984
rect 286594 2972 286600 2984
rect 280120 2944 286600 2972
rect 280120 2932 280126 2944
rect 286594 2932 286600 2944
rect 286652 2932 286658 2984
rect 404262 2932 404268 2984
rect 404320 2972 404326 2984
rect 420178 2972 420184 2984
rect 404320 2944 420184 2972
rect 404320 2932 404326 2944
rect 420178 2932 420184 2944
rect 420236 2932 420242 2984
rect 423582 2932 423588 2984
rect 423640 2972 423646 2984
rect 441522 2972 441528 2984
rect 423640 2944 441528 2972
rect 423640 2932 423646 2944
rect 441522 2932 441528 2944
rect 441580 2932 441586 2984
rect 442902 2932 442908 2984
rect 442960 2972 442966 2984
rect 442960 2944 443960 2972
rect 442960 2932 442966 2944
rect 255222 2864 255228 2916
rect 255280 2904 255286 2916
rect 259454 2904 259460 2916
rect 255280 2876 259460 2904
rect 255280 2864 255286 2876
rect 259454 2864 259460 2876
rect 259512 2864 259518 2916
rect 288342 2864 288348 2916
rect 288400 2904 288406 2916
rect 294874 2904 294880 2916
rect 288400 2876 294880 2904
rect 288400 2864 288406 2876
rect 294874 2864 294880 2876
rect 294932 2864 294938 2916
rect 426342 2864 426348 2916
rect 426400 2904 426406 2916
rect 443822 2904 443828 2916
rect 426400 2876 443828 2904
rect 426400 2864 426406 2876
rect 443822 2864 443828 2876
rect 443880 2864 443886 2916
rect 443932 2904 443960 2944
rect 447042 2932 447048 2984
rect 447100 2972 447106 2984
rect 466270 2972 466276 2984
rect 447100 2944 466276 2972
rect 447100 2932 447106 2944
rect 466270 2932 466276 2944
rect 466328 2932 466334 2984
rect 533982 2932 533988 2984
rect 534040 2972 534046 2984
rect 560846 2972 560852 2984
rect 534040 2944 560852 2972
rect 534040 2932 534046 2944
rect 560846 2932 560852 2944
rect 560904 2932 560910 2984
rect 461578 2904 461584 2916
rect 443932 2876 461584 2904
rect 461578 2864 461584 2876
rect 461636 2864 461642 2916
rect 531222 2864 531228 2916
rect 531280 2904 531286 2916
rect 557350 2904 557356 2916
rect 531280 2876 557356 2904
rect 531280 2864 531286 2876
rect 557350 2864 557356 2876
rect 557408 2864 557414 2916
rect 436002 2796 436008 2848
rect 436060 2836 436066 2848
rect 454494 2836 454500 2848
rect 436060 2808 454500 2836
rect 436060 2796 436066 2808
rect 454494 2796 454500 2808
rect 454552 2796 454558 2848
rect 454589 2839 454647 2845
rect 454589 2805 454601 2839
rect 454635 2836 454647 2839
rect 472250 2836 472256 2848
rect 454635 2808 472256 2836
rect 454635 2805 454647 2808
rect 454589 2799 454647 2805
rect 472250 2796 472256 2808
rect 472308 2796 472314 2848
rect 524322 2796 524328 2848
rect 524380 2836 524386 2848
rect 550266 2836 550272 2848
rect 524380 2808 550272 2836
rect 524380 2796 524386 2808
rect 550266 2796 550272 2808
rect 550324 2796 550330 2848
<< via1 >>
rect 154120 700952 154172 701004
rect 320180 700952 320232 701004
rect 137836 700884 137888 700936
rect 316040 700884 316092 700936
rect 246948 700816 247000 700868
rect 462320 700816 462372 700868
rect 251088 700748 251140 700800
rect 478512 700748 478564 700800
rect 89168 700680 89220 700732
rect 335360 700680 335412 700732
rect 72976 700612 73028 700664
rect 329840 700612 329892 700664
rect 331864 700612 331916 700664
rect 429844 700612 429896 700664
rect 233148 700544 233200 700596
rect 527180 700544 527232 700596
rect 40500 700476 40552 700528
rect 339500 700476 339552 700528
rect 170312 700408 170364 700460
rect 180064 700408 180116 700460
rect 237288 700408 237340 700460
rect 543464 700408 543516 700460
rect 24308 700340 24360 700392
rect 349160 700340 349212 700392
rect 8116 700272 8168 700324
rect 345020 700272 345072 700324
rect 443644 700272 443696 700324
rect 494796 700272 494848 700324
rect 266268 700204 266320 700256
rect 413652 700204 413704 700256
rect 260748 700136 260800 700188
rect 397460 700136 397512 700188
rect 202788 700068 202840 700120
rect 302240 700068 302292 700120
rect 218980 700000 219032 700052
rect 306380 700000 306432 700052
rect 280068 699932 280120 699984
rect 348792 699932 348844 699984
rect 274548 699864 274600 699916
rect 332508 699864 332560 699916
rect 235172 699796 235224 699848
rect 238024 699796 238076 699848
rect 267648 699796 267700 699848
rect 288440 699796 288492 699848
rect 283840 699728 283892 699780
rect 292580 699728 292632 699780
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 363604 699660 363656 699712
rect 364984 699660 365036 699712
rect 555424 699660 555476 699712
rect 559656 699660 559708 699712
rect 219348 696940 219400 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 353944 683204 353996 683256
rect 223488 683136 223540 683188
rect 580172 683136 580224 683188
rect 256608 676812 256660 676864
rect 331864 676812 331916 676864
rect 283932 674500 283984 674552
rect 299480 674500 299532 674552
rect 238024 674432 238076 674484
rect 298008 674432 298060 674484
rect 269856 674364 269908 674416
rect 363604 674364 363656 674416
rect 180064 674296 180116 674348
rect 312084 674296 312136 674348
rect 241704 674228 241756 674280
rect 443644 674228 443696 674280
rect 106188 674160 106240 674212
rect 326160 674160 326212 674212
rect 227536 674092 227588 674144
rect 555424 674092 555476 674144
rect 218152 673412 218204 673464
rect 219348 673412 219400 673464
rect 232320 673412 232372 673464
rect 233148 673412 233200 673464
rect 255780 673412 255832 673464
rect 256608 673412 256660 673464
rect 265164 673412 265216 673464
rect 266268 673412 266320 673464
rect 279240 673412 279292 673464
rect 280068 673412 280120 673464
rect 204352 673344 204404 673396
rect 391940 673344 391992 673396
rect 67916 673276 67968 673328
rect 359464 673276 359516 673328
rect 180616 673208 180668 673260
rect 555516 673208 555568 673260
rect 5172 673140 5224 673192
rect 406016 673140 406068 673192
rect 5080 673072 5132 673124
rect 420092 673072 420144 673124
rect 147772 673004 147824 673056
rect 566648 673004 566700 673056
rect 138388 672936 138440 672988
rect 576308 672936 576360 672988
rect 4988 672868 5040 672920
rect 448336 672868 448388 672920
rect 124312 672800 124364 672852
rect 571984 672800 572036 672852
rect 119528 672732 119580 672784
rect 572076 672732 572128 672784
rect 7840 672664 7892 672716
rect 462412 672664 462464 672716
rect 11888 672596 11940 672648
rect 476488 672596 476540 672648
rect 105452 672528 105504 672580
rect 570604 672528 570656 672580
rect 13268 672460 13320 672512
rect 490564 672460 490616 672512
rect 81992 672392 82044 672444
rect 558276 672392 558328 672444
rect 91376 672324 91428 672376
rect 573456 672324 573508 672376
rect 96068 672256 96120 672308
rect 578884 672256 578936 672308
rect 77300 672188 77352 672240
rect 569316 672188 569368 672240
rect 4804 672120 4856 672172
rect 499948 672120 500000 672172
rect 500868 672120 500920 672172
rect 542176 672120 542228 672172
rect 7748 672052 7800 672104
rect 504640 672052 504692 672104
rect 3056 671984 3108 672036
rect 363788 671984 363840 672036
rect 10692 671916 10744 671968
rect 373172 671916 373224 671968
rect 199384 671848 199436 671900
rect 565268 671848 565320 671900
rect 213460 671780 213512 671832
rect 580172 671780 580224 671832
rect 190000 671712 190052 671764
rect 556988 671712 557040 671764
rect 13452 671644 13504 671696
rect 401324 671644 401376 671696
rect 161848 671576 161900 671628
rect 554044 671576 554096 671628
rect 12072 671508 12124 671560
rect 410708 671508 410760 671560
rect 13360 671440 13412 671492
rect 424784 671440 424836 671492
rect 143080 671372 143132 671424
rect 561036 671372 561088 671424
rect 7932 671304 7984 671356
rect 438860 671304 438912 671356
rect 9036 671236 9088 671288
rect 453028 671236 453080 671288
rect 114836 671168 114888 671220
rect 565176 671168 565228 671220
rect 10416 671100 10468 671152
rect 467104 671100 467156 671152
rect 11796 671032 11848 671084
rect 481180 671032 481232 671084
rect 86684 670964 86736 671016
rect 555424 670964 555476 671016
rect 13176 670896 13228 670948
rect 495256 670896 495308 670948
rect 7656 670828 7708 670880
rect 509332 670828 509384 670880
rect 58532 670760 58584 670812
rect 573364 670760 573416 670812
rect 44456 670692 44508 670744
rect 569224 670692 569276 670744
rect 6368 670624 6420 670676
rect 359096 670624 359148 670676
rect 359464 670624 359516 670676
rect 580356 670624 580408 670676
rect 8024 670556 8076 670608
rect 368480 670556 368532 670608
rect 204076 670488 204128 670540
rect 566740 670488 566792 670540
rect 3884 670420 3936 670472
rect 204352 670420 204404 670472
rect 208768 670420 208820 670472
rect 574928 670420 574980 670472
rect 9220 670352 9272 670404
rect 377864 670352 377916 670404
rect 9128 670284 9180 670336
rect 382556 670284 382608 670336
rect 12164 670216 12216 670268
rect 387248 670216 387300 670268
rect 185308 670148 185360 670200
rect 562508 670148 562560 670200
rect 175924 670080 175976 670132
rect 555608 670080 555660 670132
rect 10600 670012 10652 670064
rect 396356 670012 396408 670064
rect 415308 670055 415360 670064
rect 415308 670021 415317 670055
rect 415317 670021 415351 670055
rect 415351 670021 415360 670055
rect 415308 670012 415360 670021
rect 433892 670012 433944 670064
rect 166816 669987 166868 669996
rect 166816 669953 166825 669987
rect 166825 669953 166859 669987
rect 166859 669953 166868 669987
rect 166816 669944 166868 669953
rect 171600 669944 171652 669996
rect 561128 669944 561180 669996
rect 157064 669876 157116 669928
rect 558368 669876 558420 669928
rect 11980 669808 12032 669860
rect 429200 669851 429252 669860
rect 429200 669817 429209 669851
rect 429209 669817 429243 669851
rect 429243 669817 429252 669851
rect 429200 669808 429252 669817
rect 443276 669851 443328 669860
rect 443276 669817 443285 669851
rect 443285 669817 443319 669851
rect 443319 669817 443328 669851
rect 443276 669808 443328 669817
rect 457444 669851 457496 669860
rect 457444 669817 457453 669851
rect 457453 669817 457487 669851
rect 457487 669817 457496 669851
rect 457444 669808 457496 669817
rect 471428 669851 471480 669860
rect 471428 669817 471437 669851
rect 471437 669817 471471 669851
rect 471471 669817 471480 669851
rect 471428 669808 471480 669817
rect 485780 669851 485832 669860
rect 485780 669817 485789 669851
rect 485789 669817 485823 669851
rect 485823 669817 485832 669851
rect 485780 669808 485832 669817
rect 500868 669851 500920 669860
rect 500868 669817 500877 669851
rect 500877 669817 500911 669851
rect 500911 669817 500920 669851
rect 500868 669808 500920 669817
rect 513748 669851 513800 669860
rect 513748 669817 513757 669851
rect 513757 669817 513791 669851
rect 513791 669817 513800 669851
rect 513748 669808 513800 669817
rect 527732 669851 527784 669860
rect 527732 669817 527741 669851
rect 527741 669817 527775 669851
rect 527775 669817 527784 669851
rect 527732 669808 527784 669817
rect 133880 669783 133932 669792
rect 133880 669749 133889 669783
rect 133889 669749 133923 669783
rect 133923 669749 133932 669783
rect 133880 669740 133932 669749
rect 152832 669740 152884 669792
rect 580448 669740 580500 669792
rect 129280 669672 129332 669724
rect 562416 669672 562468 669724
rect 110328 669604 110380 669656
rect 566556 669604 566608 669656
rect 101128 669536 101180 669588
rect 576216 669536 576268 669588
rect 63408 669511 63460 669520
rect 63408 669477 63417 669511
rect 63417 669477 63451 669511
rect 63451 669477 63460 669511
rect 63408 669468 63460 669477
rect 72976 669468 73028 669520
rect 574836 669468 574888 669520
rect 39948 669400 40000 669452
rect 560944 669400 560996 669452
rect 25964 669375 26016 669384
rect 25964 669341 25973 669375
rect 25973 669341 26007 669375
rect 26007 669341 26016 669375
rect 25964 669332 26016 669341
rect 49424 669375 49476 669384
rect 49424 669341 49433 669375
rect 49433 669341 49467 669375
rect 49467 669341 49476 669375
rect 49424 669332 49476 669341
rect 54208 669332 54260 669384
rect 580264 669332 580316 669384
rect 194692 669196 194744 669248
rect 554136 668856 554188 668908
rect 556896 668788 556948 668840
rect 6276 668720 6328 668772
rect 3792 668652 3844 668704
rect 3424 668584 3476 668636
rect 10508 668516 10560 668568
rect 578976 668448 579028 668500
rect 3700 668380 3752 668432
rect 4896 668312 4948 668364
rect 3608 668244 3660 668296
rect 3516 668176 3568 668228
rect 574744 668108 574796 668160
rect 565084 668040 565136 668092
rect 7564 667972 7616 668024
rect 562324 667904 562376 667956
rect 3240 658180 3292 658232
rect 6368 658180 6420 658232
rect 566740 644376 566792 644428
rect 580172 644376 580224 644428
rect 3332 632136 3384 632188
rect 8024 632136 8076 632188
rect 574928 632000 574980 632052
rect 579712 632000 579764 632052
rect 2964 619284 3016 619336
rect 9220 619284 9272 619336
rect 565268 618196 565320 618248
rect 579804 618196 579856 618248
rect 2872 607112 2924 607164
rect 10692 607112 10744 607164
rect 556988 591948 557040 592000
rect 580172 591948 580224 592000
rect 3148 580456 3200 580508
rect 9128 580456 9180 580508
rect 554136 578144 554188 578196
rect 580172 578144 580224 578196
rect 562508 564340 562560 564392
rect 580172 564340 580224 564392
rect 3332 554684 3384 554736
rect 12164 554684 12216 554736
rect 555608 538160 555660 538212
rect 580172 538160 580224 538212
rect 3240 528504 3292 528556
rect 10600 528504 10652 528556
rect 555516 525716 555568 525768
rect 580172 525716 580224 525768
rect 2780 515584 2832 515636
rect 5172 515584 5224 515636
rect 561128 511912 561180 511964
rect 580172 511912 580224 511964
rect 3332 502256 3384 502308
rect 13452 502256 13504 502308
rect 554044 485732 554096 485784
rect 580172 485732 580224 485784
rect 3332 476008 3384 476060
rect 12072 476008 12124 476060
rect 556896 471928 556948 471980
rect 580172 471928 580224 471980
rect 2780 463428 2832 463480
rect 5080 463428 5132 463480
rect 558368 458124 558420 458176
rect 580172 458124 580224 458176
rect 2964 449556 3016 449608
rect 6276 449556 6328 449608
rect 566648 431876 566700 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 13360 423580 13412 423632
rect 3332 411204 3384 411256
rect 11980 411204 12032 411256
rect 561036 405628 561088 405680
rect 580172 405628 580224 405680
rect 3332 371560 3384 371612
rect 7932 371560 7984 371612
rect 576308 365644 576360 365696
rect 579988 365644 580040 365696
rect 2780 358436 2832 358488
rect 4988 358436 5040 358488
rect 562416 353200 562468 353252
rect 580172 353200 580224 353252
rect 2964 346332 3016 346384
rect 10508 346332 10560 346384
rect 572076 325592 572128 325644
rect 580172 325592 580224 325644
rect 3240 320016 3292 320068
rect 9036 320016 9088 320068
rect 571984 313216 572036 313268
rect 580172 313216 580224 313268
rect 3332 306212 3384 306264
rect 7840 306212 7892 306264
rect 565176 299412 565228 299464
rect 580172 299412 580224 299464
rect 570604 273164 570656 273216
rect 580172 273164 580224 273216
rect 3240 267656 3292 267708
rect 10416 267656 10468 267708
rect 566556 259360 566608 259412
rect 579620 259360 579672 259412
rect 3332 255212 3384 255264
rect 11888 255212 11940 255264
rect 576216 245556 576268 245608
rect 580172 245556 580224 245608
rect 2780 241068 2832 241120
rect 4896 241068 4948 241120
rect 573456 233180 573508 233232
rect 580172 233180 580224 233232
rect 3332 215228 3384 215280
rect 11796 215228 11848 215280
rect 555424 206932 555476 206984
rect 579896 206932 579948 206984
rect 3332 202784 3384 202836
rect 13268 202784 13320 202836
rect 569316 193128 569368 193180
rect 580172 193128 580224 193180
rect 558276 179324 558328 179376
rect 580172 179324 580224 179376
rect 574836 166948 574888 167000
rect 580172 166948 580224 167000
rect 3332 164160 3384 164212
rect 13176 164160 13228 164212
rect 574744 153144 574796 153196
rect 579620 153144 579672 153196
rect 3608 150356 3660 150408
rect 7748 150356 7800 150408
rect 2780 136824 2832 136876
rect 4804 136824 4856 136876
rect 573364 126896 573416 126948
rect 580172 126896 580224 126948
rect 565084 113092 565136 113144
rect 580172 113092 580224 113144
rect 2964 111120 3016 111172
rect 7656 111120 7708 111172
rect 3240 97928 3292 97980
rect 11704 97928 11756 97980
rect 569224 86912 569276 86964
rect 580172 86912 580224 86964
rect 576124 73108 576176 73160
rect 580172 73108 580224 73160
rect 3516 71612 3568 71664
rect 8944 71612 8996 71664
rect 560944 60664 560996 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 13084 59304 13136 59356
rect 171140 48288 171192 48340
rect 12256 48220 12308 48272
rect 24308 48220 24360 48272
rect 27436 48220 27488 48272
rect 38476 48220 38528 48272
rect 45468 48220 45520 48272
rect 54944 48220 54996 48272
rect 172152 48220 172204 48272
rect 4068 48152 4120 48204
rect 16580 48152 16632 48204
rect 17868 48152 17920 48204
rect 29736 48152 29788 48204
rect 33048 48152 33100 48204
rect 43996 48152 44048 48204
rect 48228 48152 48280 48204
rect 58256 48152 58308 48204
rect 59268 48152 59320 48204
rect 68100 48152 68152 48204
rect 73068 48152 73120 48204
rect 81256 48152 81308 48204
rect 8208 48084 8260 48136
rect 20996 48084 21048 48136
rect 24768 48084 24820 48136
rect 36360 48084 36412 48136
rect 41328 48084 41380 48136
rect 51632 48084 51684 48136
rect 52368 48084 52420 48136
rect 61476 48084 61528 48136
rect 67548 48084 67600 48136
rect 75736 48084 75788 48136
rect 95056 48084 95108 48136
rect 102048 48084 102100 48136
rect 12348 48016 12400 48068
rect 25412 48016 25464 48068
rect 28908 48016 28960 48068
rect 39580 48016 39632 48068
rect 39948 48016 40000 48068
rect 50528 48016 50580 48068
rect 50988 48016 51040 48068
rect 60464 48016 60516 48068
rect 61936 48016 61988 48068
rect 70308 48016 70360 48068
rect 13728 47948 13780 48000
rect 26424 47948 26476 48000
rect 30288 47948 30340 48000
rect 41788 47948 41840 48000
rect 42708 47948 42760 48000
rect 52736 47948 52788 48000
rect 62028 47948 62080 48000
rect 71412 47948 71464 48000
rect 6828 47880 6880 47932
rect 19892 47880 19944 47932
rect 26148 47880 26200 47932
rect 37464 47880 37516 47932
rect 38568 47880 38620 47932
rect 49516 47880 49568 47932
rect 53656 47880 53708 47932
rect 62580 47880 62632 47932
rect 63408 47880 63460 47932
rect 5448 47812 5500 47864
rect 18788 47812 18840 47864
rect 19248 47812 19300 47864
rect 30840 47812 30892 47864
rect 31668 47812 31720 47864
rect 42892 47812 42944 47864
rect 44088 47812 44140 47864
rect 53840 47812 53892 47864
rect 55128 47812 55180 47864
rect 64788 47812 64840 47864
rect 70308 47880 70360 47932
rect 77944 48016 77996 48068
rect 79968 48016 80020 48068
rect 87788 48016 87840 48068
rect 91008 48016 91060 48068
rect 97632 48016 97684 48068
rect 92388 47948 92440 48000
rect 98736 47948 98788 48000
rect 102048 47948 102100 48000
rect 107568 47948 107620 48000
rect 531412 47948 531464 48000
rect 74448 47880 74500 47932
rect 82360 47880 82412 47932
rect 86776 47880 86828 47932
rect 93308 47880 93360 47932
rect 103336 47880 103388 47932
rect 108580 47880 108632 47932
rect 115848 47880 115900 47932
rect 120632 47880 120684 47932
rect 135168 47880 135220 47932
rect 138204 47880 138256 47932
rect 146208 47880 146260 47932
rect 149152 47880 149204 47932
rect 158628 47880 158680 47932
rect 160100 47880 160152 47932
rect 212724 47880 212776 47932
rect 214012 47880 214064 47932
rect 536932 47948 536984 48000
rect 538128 47948 538180 48000
rect 546776 47948 546828 48000
rect 547788 47948 547840 48000
rect 547880 47948 547932 48000
rect 549076 47948 549128 48000
rect 557540 47880 557592 47932
rect 72516 47812 72568 47864
rect 2688 47744 2740 47796
rect 15476 47744 15528 47796
rect 20628 47744 20680 47796
rect 31944 47744 31996 47796
rect 35808 47744 35860 47796
rect 46204 47744 46256 47796
rect 46848 47744 46900 47796
rect 57152 47744 57204 47796
rect 57888 47744 57940 47796
rect 66996 47744 67048 47796
rect 9588 47676 9640 47728
rect 22100 47676 22152 47728
rect 23388 47676 23440 47728
rect 35256 47676 35308 47728
rect 37096 47676 37148 47728
rect 47308 47676 47360 47728
rect 53748 47676 53800 47728
rect 63684 47676 63736 47728
rect 64788 47676 64840 47728
rect 3976 47608 4028 47660
rect 17684 47608 17736 47660
rect 28816 47608 28868 47660
rect 40684 47608 40736 47660
rect 45376 47608 45428 47660
rect 56048 47608 56100 47660
rect 56508 47608 56560 47660
rect 65892 47608 65944 47660
rect 66168 47676 66220 47728
rect 74632 47812 74684 47864
rect 84108 47812 84160 47864
rect 91100 47812 91152 47864
rect 93768 47812 93820 47864
rect 99840 47812 99892 47864
rect 107568 47812 107620 47864
rect 112996 47812 113048 47864
rect 114468 47812 114520 47864
rect 119620 47812 119672 47864
rect 130384 47812 130436 47864
rect 131672 47812 131724 47864
rect 137284 47812 137336 47864
rect 140412 47812 140464 47864
rect 144828 47812 144880 47864
rect 146944 47812 146996 47864
rect 148968 47812 149020 47864
rect 151360 47812 151412 47864
rect 153108 47812 153160 47864
rect 154672 47812 154724 47864
rect 155868 47812 155920 47864
rect 157892 47812 157944 47864
rect 160008 47812 160060 47864
rect 161204 47812 161256 47864
rect 162768 47812 162820 47864
rect 164516 47812 164568 47864
rect 166908 47812 166960 47864
rect 167736 47812 167788 47864
rect 176660 47812 176712 47864
rect 177672 47812 177724 47864
rect 186320 47812 186372 47864
rect 187516 47812 187568 47864
rect 206100 47812 206152 47864
rect 206928 47812 206980 47864
rect 217048 47812 217100 47864
rect 217968 47812 218020 47864
rect 222568 47812 222620 47864
rect 223488 47812 223540 47864
rect 226892 47812 226944 47864
rect 227628 47812 227680 47864
rect 227996 47812 228048 47864
rect 229008 47812 229060 47864
rect 229100 47812 229152 47864
rect 231952 47812 232004 47864
rect 232412 47812 232464 47864
rect 233148 47812 233200 47864
rect 233516 47812 233568 47864
rect 234528 47812 234580 47864
rect 234620 47812 234672 47864
rect 237472 47812 237524 47864
rect 237840 47812 237892 47864
rect 238668 47812 238720 47864
rect 240048 47812 240100 47864
rect 240784 47812 240836 47864
rect 244464 47812 244516 47864
rect 245568 47812 245620 47864
rect 248880 47812 248932 47864
rect 249708 47812 249760 47864
rect 249892 47812 249944 47864
rect 250996 47812 251048 47864
rect 254308 47812 254360 47864
rect 255228 47812 255280 47864
rect 255412 47812 255464 47864
rect 256516 47812 256568 47864
rect 260932 47812 260984 47864
rect 264244 47812 264296 47864
rect 270776 47812 270828 47864
rect 271788 47812 271840 47864
rect 281724 47812 281776 47864
rect 282736 47812 282788 47864
rect 286048 47812 286100 47864
rect 286968 47812 287020 47864
rect 287152 47812 287204 47864
rect 288348 47812 288400 47864
rect 291568 47812 291620 47864
rect 292488 47812 292540 47864
rect 292672 47812 292724 47864
rect 293776 47812 293828 47864
rect 296996 47812 297048 47864
rect 298008 47812 298060 47864
rect 301412 47812 301464 47864
rect 302148 47812 302200 47864
rect 302516 47812 302568 47864
rect 303528 47812 303580 47864
rect 303620 47812 303672 47864
rect 304908 47812 304960 47864
rect 307944 47812 307996 47864
rect 308956 47812 309008 47864
rect 312360 47812 312412 47864
rect 313188 47812 313240 47864
rect 317880 47812 317932 47864
rect 318708 47812 318760 47864
rect 324412 47812 324464 47864
rect 325516 47812 325568 47864
rect 328828 47812 328880 47864
rect 329748 47812 329800 47864
rect 329932 47812 329984 47864
rect 331128 47812 331180 47864
rect 334256 47812 334308 47864
rect 335268 47812 335320 47864
rect 335360 47812 335412 47864
rect 336648 47812 336700 47864
rect 339776 47812 339828 47864
rect 340788 47812 340840 47864
rect 350724 47812 350776 47864
rect 351736 47812 351788 47864
rect 355048 47812 355100 47864
rect 355968 47812 356020 47864
rect 360568 47812 360620 47864
rect 361488 47812 361540 47864
rect 366088 47812 366140 47864
rect 367008 47812 367060 47864
rect 367100 47812 367152 47864
rect 368296 47812 368348 47864
rect 371516 47812 371568 47864
rect 372528 47812 372580 47864
rect 372620 47812 372672 47864
rect 373816 47812 373868 47864
rect 375932 47812 375984 47864
rect 376668 47812 376720 47864
rect 377036 47812 377088 47864
rect 378048 47812 378100 47864
rect 378140 47812 378192 47864
rect 379428 47812 379480 47864
rect 382464 47812 382516 47864
rect 383476 47812 383528 47864
rect 386880 47812 386932 47864
rect 387708 47812 387760 47864
rect 387984 47812 388036 47864
rect 389088 47812 389140 47864
rect 392308 47812 392360 47864
rect 393228 47812 393280 47864
rect 403256 47812 403308 47864
rect 404268 47812 404320 47864
rect 404360 47812 404412 47864
rect 405648 47812 405700 47864
rect 408776 47812 408828 47864
rect 409788 47812 409840 47864
rect 409880 47812 409932 47864
rect 411076 47812 411128 47864
rect 418620 47812 418672 47864
rect 419448 47812 419500 47864
rect 419724 47812 419776 47864
rect 420736 47812 420788 47864
rect 429568 47812 429620 47864
rect 430488 47812 430540 47864
rect 430672 47812 430724 47864
rect 431868 47812 431920 47864
rect 436192 47812 436244 47864
rect 437296 47812 437348 47864
rect 439412 47812 439464 47864
rect 440148 47812 440200 47864
rect 440516 47812 440568 47864
rect 441528 47812 441580 47864
rect 441620 47812 441672 47864
rect 442908 47812 442960 47864
rect 446036 47812 446088 47864
rect 447048 47812 447100 47864
rect 450360 47812 450412 47864
rect 451188 47812 451240 47864
rect 451464 47812 451516 47864
rect 452568 47812 452620 47864
rect 456984 47812 457036 47864
rect 457996 47812 458048 47864
rect 461308 47812 461360 47864
rect 462228 47812 462280 47864
rect 466828 47812 466880 47864
rect 467748 47812 467800 47864
rect 467932 47812 467984 47864
rect 469128 47812 469180 47864
rect 472256 47812 472308 47864
rect 473268 47812 473320 47864
rect 473360 47812 473412 47864
rect 474556 47812 474608 47864
rect 477776 47812 477828 47864
rect 478788 47812 478840 47864
rect 478880 47812 478932 47864
rect 480076 47812 480128 47864
rect 483296 47812 483348 47864
rect 484216 47812 484268 47864
rect 493140 47812 493192 47864
rect 493968 47812 494020 47864
rect 494244 47812 494296 47864
rect 495348 47812 495400 47864
rect 499672 47812 499724 47864
rect 500776 47812 500828 47864
rect 504088 47812 504140 47864
rect 505008 47812 505060 47864
rect 508412 47812 508464 47864
rect 509148 47812 509200 47864
rect 510620 47812 510672 47864
rect 511908 47812 511960 47864
rect 513932 47812 513984 47864
rect 514668 47812 514720 47864
rect 515036 47812 515088 47864
rect 516048 47812 516100 47864
rect 516140 47812 516192 47864
rect 517428 47812 517480 47864
rect 519360 47812 519412 47864
rect 520188 47812 520240 47864
rect 520464 47812 520516 47864
rect 521568 47812 521620 47864
rect 524880 47812 524932 47864
rect 525708 47812 525760 47864
rect 525984 47812 526036 47864
rect 526996 47812 527048 47864
rect 530400 47812 530452 47864
rect 531228 47812 531280 47864
rect 535828 47812 535880 47864
rect 536748 47812 536800 47864
rect 77208 47744 77260 47796
rect 84568 47744 84620 47796
rect 86868 47744 86920 47796
rect 94412 47744 94464 47796
rect 100668 47744 100720 47796
rect 106464 47744 106516 47796
rect 113088 47744 113140 47796
rect 118516 47744 118568 47796
rect 121368 47744 121420 47796
rect 126152 47744 126204 47796
rect 126888 47744 126940 47796
rect 130568 47744 130620 47796
rect 132408 47744 132460 47796
rect 135996 47744 136048 47796
rect 136548 47744 136600 47796
rect 139308 47744 139360 47796
rect 147588 47744 147640 47796
rect 150256 47744 150308 47796
rect 153016 47744 153068 47796
rect 155684 47744 155736 47796
rect 193312 47744 193364 47796
rect 194048 47744 194100 47796
rect 211620 47744 211672 47796
rect 212724 47744 212776 47796
rect 225788 47744 225840 47796
rect 227812 47744 227864 47796
rect 243360 47744 243412 47796
rect 246304 47744 246356 47796
rect 306932 47744 306984 47796
rect 307668 47744 307720 47796
rect 318984 47744 319036 47796
rect 320088 47744 320140 47796
rect 370412 47744 370464 47796
rect 371148 47744 371200 47796
rect 435088 47744 435140 47796
rect 436008 47744 436060 47796
rect 534724 47744 534776 47796
rect 560944 47812 560996 47864
rect 538036 47744 538088 47796
rect 564532 47744 564584 47796
rect 85488 47676 85540 47728
rect 92204 47676 92256 47728
rect 103428 47676 103480 47728
rect 109684 47676 109736 47728
rect 111616 47676 111668 47728
rect 116308 47676 116360 47728
rect 117228 47676 117280 47728
rect 121736 47676 121788 47728
rect 122748 47676 122800 47728
rect 127256 47676 127308 47728
rect 137928 47676 137980 47728
rect 141516 47676 141568 47728
rect 238944 47676 238996 47728
rect 240048 47676 240100 47728
rect 340880 47676 340932 47728
rect 342076 47676 342128 47728
rect 498568 47676 498620 47728
rect 502984 47676 503036 47728
rect 509516 47676 509568 47728
rect 510528 47676 510580 47728
rect 528192 47676 528244 47728
rect 552296 47676 552348 47728
rect 553308 47676 553360 47728
rect 1308 47540 1360 47592
rect 14464 47540 14516 47592
rect 20536 47540 20588 47592
rect 32772 47540 32824 47592
rect 37188 47540 37240 47592
rect 48412 47540 48464 47592
rect 49608 47540 49660 47592
rect 59360 47540 59412 47592
rect 60648 47540 60700 47592
rect 69204 47540 69256 47592
rect 10968 47472 11020 47524
rect 23204 47472 23256 47524
rect 34428 47472 34480 47524
rect 45100 47472 45152 47524
rect 71688 47608 71740 47660
rect 80152 47608 80204 47660
rect 81348 47608 81400 47660
rect 88892 47608 88944 47660
rect 89628 47608 89680 47660
rect 96620 47608 96672 47660
rect 104808 47608 104860 47660
rect 110788 47608 110840 47660
rect 111708 47608 111760 47660
rect 117412 47608 117464 47660
rect 157248 47608 157300 47660
rect 158996 47608 159048 47660
rect 164148 47608 164200 47660
rect 165620 47608 165672 47660
rect 218152 47608 218204 47660
rect 219348 47608 219400 47660
rect 221464 47608 221516 47660
rect 222844 47608 222896 47660
rect 223672 47608 223724 47660
rect 224776 47608 224828 47660
rect 266360 47608 266412 47660
rect 267648 47608 267700 47660
rect 276204 47608 276256 47660
rect 277308 47608 277360 47660
rect 313464 47608 313516 47660
rect 314568 47608 314620 47660
rect 356152 47608 356204 47660
rect 357348 47608 357400 47660
rect 361672 47608 361724 47660
rect 362868 47608 362920 47660
rect 495256 47608 495308 47660
rect 504364 47608 504416 47660
rect 505192 47608 505244 47660
rect 515404 47608 515456 47660
rect 541348 47608 541400 47660
rect 568580 47608 568632 47660
rect 70216 47540 70268 47592
rect 79048 47540 79100 47592
rect 82728 47540 82780 47592
rect 89996 47540 90048 47592
rect 106188 47540 106240 47592
rect 111892 47540 111944 47592
rect 259828 47540 259880 47592
rect 260748 47540 260800 47592
rect 265256 47540 265308 47592
rect 270592 47540 270644 47592
rect 275100 47540 275152 47592
rect 275928 47540 275980 47592
rect 280620 47540 280672 47592
rect 281448 47540 281500 47592
rect 323308 47540 323360 47592
rect 324228 47540 324280 47592
rect 344100 47540 344152 47592
rect 344928 47540 344980 47592
rect 349620 47540 349672 47592
rect 350448 47540 350500 47592
rect 381360 47540 381412 47592
rect 382188 47540 382240 47592
rect 397828 47540 397880 47592
rect 398748 47540 398800 47592
rect 424140 47540 424192 47592
rect 424968 47540 425020 47592
rect 444932 47540 444984 47592
rect 445668 47540 445720 47592
rect 455880 47540 455932 47592
rect 456708 47540 456760 47592
rect 462412 47540 462464 47592
rect 482284 47540 482336 47592
rect 487620 47540 487672 47592
rect 488448 47540 488500 47592
rect 488724 47540 488776 47592
rect 512092 47540 512144 47592
rect 553400 47540 553452 47592
rect 73528 47472 73580 47524
rect 393412 47472 393464 47524
rect 394516 47472 394568 47524
rect 554780 47472 554832 47524
rect 15108 47404 15160 47456
rect 27528 47404 27580 47456
rect 75828 47404 75880 47456
rect 83464 47404 83516 47456
rect 96528 47404 96580 47456
rect 103152 47404 103204 47456
rect 143448 47404 143500 47456
rect 145840 47404 145892 47456
rect 345204 47404 345256 47456
rect 346308 47404 346360 47456
rect 398932 47404 398984 47456
rect 400036 47404 400088 47456
rect 414204 47404 414256 47456
rect 415308 47404 415360 47456
rect 425244 47404 425296 47456
rect 426348 47404 426400 47456
rect 447140 47404 447192 47456
rect 448428 47404 448480 47456
rect 16488 47336 16540 47388
rect 28632 47336 28684 47388
rect 22008 47268 22060 47320
rect 34152 47268 34204 47320
rect 95148 47268 95200 47320
rect 100944 47268 100996 47320
rect 124128 47268 124180 47320
rect 128360 47268 128412 47320
rect 207204 47268 207256 47320
rect 208492 47268 208544 47320
rect 298100 47268 298152 47320
rect 299296 47268 299348 47320
rect 492036 47268 492088 47320
rect 497464 47268 497516 47320
rect 542452 47268 542504 47320
rect 543648 47268 543700 47320
rect 119896 47132 119948 47184
rect 125048 47132 125100 47184
rect 128268 47132 128320 47184
rect 132684 47132 132736 47184
rect 110328 47064 110380 47116
rect 115204 47064 115256 47116
rect 131028 47064 131080 47116
rect 134892 47064 134944 47116
rect 139308 47064 139360 47116
rect 142620 47064 142672 47116
rect 78496 46996 78548 47048
rect 86684 46996 86736 47048
rect 99288 46996 99340 47048
rect 105360 46996 105412 47048
rect 108948 46996 109000 47048
rect 114100 46996 114152 47048
rect 118608 46996 118660 47048
rect 122840 46996 122892 47048
rect 125508 46996 125560 47048
rect 129464 46996 129516 47048
rect 129648 46996 129700 47048
rect 133788 46996 133840 47048
rect 140688 46996 140740 47048
rect 143632 46996 143684 47048
rect 151728 46996 151780 47048
rect 153568 46996 153620 47048
rect 271880 46996 271932 47048
rect 277492 46996 277544 47048
rect 68928 46928 68980 46980
rect 76840 46928 76892 46980
rect 78588 46928 78640 46980
rect 85580 46928 85632 46980
rect 88248 46928 88300 46980
rect 95516 46928 95568 46980
rect 97908 46928 97960 46980
rect 104256 46928 104308 46980
rect 119988 46928 120040 46980
rect 123944 46928 123996 46980
rect 137100 46928 137152 46980
rect 142068 46928 142120 46980
rect 144736 46928 144788 46980
rect 133788 46860 133840 46912
rect 148048 46928 148100 46980
rect 151084 46928 151136 46980
rect 152464 46928 152516 46980
rect 161296 46928 161348 46980
rect 163412 46928 163464 46980
rect 199568 46928 199620 46980
rect 200212 46928 200264 46980
rect 219256 46928 219308 46980
rect 220084 46928 220136 46980
rect 566464 46860 566516 46912
rect 580172 46860 580224 46912
rect 144828 46724 144880 46776
rect 3516 45500 3568 45552
rect 7564 45500 7616 45552
rect 558184 33056 558236 33108
rect 580172 33056 580224 33108
rect 2780 32920 2832 32972
rect 6184 32920 6236 32972
rect 3516 20612 3568 20664
rect 10324 20612 10376 20664
rect 562324 20612 562376 20664
rect 579988 20612 580040 20664
rect 474556 11840 474608 11892
rect 474648 11636 474700 11688
rect 515404 7692 515456 7744
rect 530124 7692 530176 7744
rect 480076 7624 480128 7676
rect 501788 7624 501840 7676
rect 504364 7624 504416 7676
rect 519544 7624 519596 7676
rect 469036 7556 469088 7608
rect 491116 7556 491168 7608
rect 497464 7556 497516 7608
rect 515956 7556 516008 7608
rect 516048 7556 516100 7608
rect 540796 7556 540848 7608
rect 556804 6808 556856 6860
rect 580172 6808 580224 6860
rect 560944 5516 560996 5568
rect 562048 5516 562100 5568
rect 502984 5176 503036 5228
rect 523040 5176 523092 5228
rect 509148 5108 509200 5160
rect 533712 5108 533764 5160
rect 473268 5040 473320 5092
rect 494704 5040 494756 5092
rect 502248 5040 502300 5092
rect 526628 5040 526680 5092
rect 466368 4972 466420 5024
rect 487620 4972 487672 5024
rect 518808 4972 518860 5024
rect 544384 4972 544436 5024
rect 485688 4904 485740 4956
rect 508872 4904 508924 4956
rect 525708 4904 525760 4956
rect 551468 4904 551520 4956
rect 476028 4836 476080 4888
rect 498200 4836 498252 4888
rect 511816 4836 511868 4888
rect 537208 4836 537260 4888
rect 459468 4768 459520 4820
rect 480536 4768 480588 4820
rect 482928 4768 482980 4820
rect 505376 4768 505428 4820
rect 521476 4768 521528 4820
rect 547880 4768 547932 4820
rect 482284 4156 482336 4208
rect 484032 4156 484084 4208
rect 209688 4088 209740 4140
rect 210976 4088 211028 4140
rect 229008 4088 229060 4140
rect 231032 4088 231084 4140
rect 237288 4088 237340 4140
rect 240508 4088 240560 4140
rect 256516 4088 256568 4140
rect 260656 4088 260708 4140
rect 262128 4088 262180 4140
rect 267740 4088 267792 4140
rect 282736 4088 282788 4140
rect 288992 4088 289044 4140
rect 253848 4020 253900 4072
rect 258264 4020 258316 4072
rect 304908 4020 304960 4072
rect 312636 4020 312688 4072
rect 314568 4020 314620 4072
rect 323308 4088 323360 4140
rect 324228 4088 324280 4140
rect 333888 4088 333940 4140
rect 343548 4088 343600 4140
rect 355232 4088 355284 4140
rect 355968 4088 356020 4140
rect 368204 4088 368256 4140
rect 371148 4088 371200 4140
rect 384764 4088 384816 4140
rect 384948 4088 385000 4140
rect 399944 4088 399996 4140
rect 411076 4088 411128 4140
rect 427268 4088 427320 4140
rect 429108 4088 429160 4140
rect 447416 4088 447468 4140
rect 451188 4088 451240 4140
rect 471060 4088 471112 4140
rect 477408 4088 477460 4140
rect 499396 4088 499448 4140
rect 505008 4088 505060 4140
rect 529020 4088 529072 4140
rect 529848 4088 529900 4140
rect 556160 4088 556212 4140
rect 245476 3952 245528 4004
rect 249984 3952 250036 4004
rect 264888 3952 264940 4004
rect 270040 3952 270092 4004
rect 281448 3952 281500 4004
rect 287796 3952 287848 4004
rect 293776 3952 293828 4004
rect 300768 3952 300820 4004
rect 311808 3952 311860 4004
rect 320916 4020 320968 4072
rect 331128 4020 331180 4072
rect 340972 4020 341024 4072
rect 342076 4020 342128 4072
rect 352840 4020 352892 4072
rect 354588 4020 354640 4072
rect 366916 4020 366968 4072
rect 373816 4020 373868 4072
rect 387156 4020 387208 4072
rect 394516 4020 394568 4072
rect 409604 4020 409656 4072
rect 416688 4020 416740 4072
rect 434444 4020 434496 4072
rect 434628 4020 434680 4072
rect 453304 4020 453356 4072
rect 456708 4020 456760 4072
rect 476948 4020 477000 4072
rect 481548 4020 481600 4072
rect 504180 4020 504232 4072
rect 510528 4020 510580 4072
rect 534908 4020 534960 4072
rect 543648 4020 543700 4072
rect 570328 4020 570380 4072
rect 317328 3952 317380 4004
rect 332508 3952 332560 4004
rect 343364 3952 343416 4004
rect 346308 3952 346360 4004
rect 357532 3952 357584 4004
rect 365628 3952 365680 4004
rect 378876 3952 378928 4004
rect 382188 3952 382240 4004
rect 396540 3952 396592 4004
rect 398748 3952 398800 4004
rect 414296 3952 414348 4004
rect 420736 3952 420788 4004
rect 437940 3952 437992 4004
rect 441528 3952 441580 4004
rect 460388 3952 460440 4004
rect 463608 3952 463660 4004
rect 485228 3952 485280 4004
rect 487068 3952 487120 4004
rect 510068 3952 510120 4004
rect 514668 3952 514720 4004
rect 539600 3952 539652 4004
rect 546408 3952 546460 4004
rect 573916 3952 573968 4004
rect 303528 3884 303580 3936
rect 311440 3884 311492 3936
rect 326804 3884 326856 3936
rect 326988 3884 327040 3936
rect 337476 3884 337528 3936
rect 342168 3884 342220 3936
rect 354036 3884 354088 3936
rect 248328 3816 248380 3868
rect 252376 3816 252428 3868
rect 274548 3816 274600 3868
rect 280712 3816 280764 3868
rect 292488 3816 292540 3868
rect 299664 3816 299716 3868
rect 308956 3816 309008 3868
rect 317328 3816 317380 3868
rect 318708 3816 318760 3868
rect 328000 3816 328052 3868
rect 328368 3816 328420 3868
rect 338672 3816 338724 3868
rect 339408 3816 339460 3868
rect 350448 3816 350500 3868
rect 351736 3816 351788 3868
rect 286968 3748 287020 3800
rect 293684 3748 293736 3800
rect 309048 3748 309100 3800
rect 318524 3748 318576 3800
rect 320088 3748 320140 3800
rect 329196 3748 329248 3800
rect 329748 3748 329800 3800
rect 339868 3748 339920 3800
rect 347688 3748 347740 3800
rect 359924 3816 359976 3868
rect 360108 3884 360160 3936
rect 372896 3884 372948 3936
rect 373908 3884 373960 3936
rect 388260 3884 388312 3936
rect 394608 3884 394660 3936
rect 410800 3884 410852 3936
rect 412548 3884 412600 3936
rect 429660 3884 429712 3936
rect 430488 3884 430540 3936
rect 448612 3884 448664 3936
rect 457996 3884 458048 3936
rect 478144 3884 478196 3936
rect 484308 3884 484360 3936
rect 507676 3884 507728 3936
rect 507768 3884 507820 3936
rect 532516 3884 532568 3936
rect 539508 3884 539560 3936
rect 566832 3884 566884 3936
rect 363512 3816 363564 3868
rect 367008 3816 367060 3868
rect 379980 3816 380032 3868
rect 383476 3816 383528 3868
rect 397736 3816 397788 3868
rect 400128 3816 400180 3868
rect 416688 3816 416740 3868
rect 422208 3816 422260 3868
rect 440332 3816 440384 3868
rect 444288 3816 444340 3868
rect 463976 3816 464028 3868
rect 470508 3816 470560 3868
rect 492312 3816 492364 3868
rect 493968 3816 494020 3868
rect 517152 3816 517204 3868
rect 521568 3816 521620 3868
rect 546684 3816 546736 3868
rect 549076 3816 549128 3868
rect 576308 3816 576360 3868
rect 358728 3748 358780 3800
rect 235908 3680 235960 3732
rect 239312 3680 239364 3732
rect 267648 3680 267700 3732
rect 272432 3680 272484 3732
rect 275928 3680 275980 3732
rect 281908 3680 281960 3732
rect 284208 3680 284260 3732
rect 291384 3680 291436 3732
rect 295248 3680 295300 3732
rect 303160 3680 303212 3732
rect 306288 3680 306340 3732
rect 315028 3680 315080 3732
rect 315948 3680 316000 3732
rect 238668 3612 238720 3664
rect 241704 3612 241756 3664
rect 257988 3612 258040 3664
rect 262956 3612 263008 3664
rect 277308 3612 277360 3664
rect 283104 3612 283156 3664
rect 285588 3612 285640 3664
rect 292580 3612 292632 3664
rect 293868 3612 293920 3664
rect 301964 3612 302016 3664
rect 302148 3612 302200 3664
rect 310244 3612 310296 3664
rect 313188 3612 313240 3664
rect 322112 3612 322164 3664
rect 325516 3680 325568 3732
rect 335084 3680 335136 3732
rect 336648 3680 336700 3732
rect 346952 3680 347004 3732
rect 349068 3680 349120 3732
rect 325608 3612 325660 3664
rect 331036 3612 331088 3664
rect 2872 3544 2924 3596
rect 3976 3544 4028 3596
rect 19432 3544 19484 3596
rect 20536 3544 20588 3596
rect 27712 3544 27764 3596
rect 28816 3544 28868 3596
rect 44272 3544 44324 3596
rect 45376 3544 45428 3596
rect 69112 3544 69164 3596
rect 70216 3544 70268 3596
rect 77392 3544 77444 3596
rect 78496 3544 78548 3596
rect 93952 3544 94004 3596
rect 95056 3544 95108 3596
rect 168380 3544 168432 3596
rect 169668 3544 169720 3596
rect 186320 3544 186372 3596
rect 187332 3544 187384 3596
rect 201500 3544 201552 3596
rect 202696 3544 202748 3596
rect 219348 3544 219400 3596
rect 220452 3544 220504 3596
rect 223488 3544 223540 3596
rect 225144 3544 225196 3596
rect 242808 3544 242860 3596
rect 246396 3544 246448 3596
rect 251088 3544 251140 3596
rect 255872 3544 255924 3596
rect 282828 3544 282880 3596
rect 290188 3544 290240 3596
rect 299388 3544 299440 3596
rect 307944 3544 307996 3596
rect 310428 3544 310480 3596
rect 319720 3544 319772 3596
rect 322848 3544 322900 3596
rect 332692 3544 332744 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12256 3476 12308 3528
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 35992 3476 36044 3528
rect 37096 3476 37148 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 51356 3476 51408 3528
rect 52368 3476 52420 3528
rect 52552 3476 52604 3528
rect 53656 3476 53708 3528
rect 56048 3476 56100 3528
rect 56508 3476 56560 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 60832 3476 60884 3528
rect 61936 3476 61988 3528
rect 64328 3476 64380 3528
rect 64788 3476 64840 3528
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 66720 3476 66772 3528
rect 67548 3476 67600 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 82084 3476 82136 3528
rect 82728 3476 82780 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 92388 3476 92440 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 101036 3476 101088 3528
rect 102048 3476 102100 3528
rect 102232 3476 102284 3528
rect 103244 3476 103296 3528
rect 105728 3476 105780 3528
rect 106188 3476 106240 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 109316 3476 109368 3528
rect 110328 3476 110380 3528
rect 110512 3476 110564 3528
rect 111524 3476 111576 3528
rect 114008 3476 114060 3528
rect 114468 3476 114520 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 116400 3476 116452 3528
rect 117228 3476 117280 3528
rect 117596 3476 117648 3528
rect 118608 3476 118660 3528
rect 118792 3476 118844 3528
rect 119988 3476 120040 3528
rect 122288 3476 122340 3528
rect 122748 3476 122800 3528
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 125876 3476 125928 3528
rect 126888 3476 126940 3528
rect 130568 3476 130620 3528
rect 131028 3476 131080 3528
rect 132960 3476 133012 3528
rect 133788 3476 133840 3528
rect 134156 3476 134208 3528
rect 135168 3476 135220 3528
rect 136456 3476 136508 3528
rect 137284 3476 137336 3528
rect 138848 3476 138900 3528
rect 139308 3476 139360 3528
rect 140044 3476 140096 3528
rect 140688 3476 140740 3528
rect 141240 3476 141292 3528
rect 142068 3476 142120 3528
rect 142436 3476 142488 3528
rect 143448 3476 143500 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 148324 3476 148376 3528
rect 148968 3476 149020 3528
rect 149520 3476 149572 3528
rect 151084 3476 151136 3528
rect 151820 3476 151872 3528
rect 153108 3476 153160 3528
rect 154212 3476 154264 3528
rect 156052 3476 156104 3528
rect 156604 3476 156656 3528
rect 157248 3476 157300 3528
rect 157800 3476 157852 3528
rect 158628 3476 158680 3528
rect 158904 3476 158956 3528
rect 160008 3476 160060 3528
rect 160100 3476 160152 3528
rect 161388 3476 161440 3528
rect 163688 3476 163740 3528
rect 164148 3476 164200 3528
rect 164884 3476 164936 3528
rect 165712 3476 165764 3528
rect 166080 3476 166132 3528
rect 166908 3476 166960 3528
rect 167184 3476 167236 3528
rect 168564 3476 168616 3528
rect 171968 3476 172020 3528
rect 172612 3476 172664 3528
rect 173164 3476 173216 3528
rect 173808 3476 173860 3528
rect 174268 3476 174320 3528
rect 175188 3476 175240 3528
rect 179052 3476 179104 3528
rect 179512 3476 179564 3528
rect 180248 3476 180300 3528
rect 180708 3476 180760 3528
rect 180984 3476 181036 3528
rect 181444 3476 181496 3528
rect 187700 3476 187752 3528
rect 188528 3476 188580 3528
rect 189080 3476 189132 3528
rect 189724 3476 189776 3528
rect 194600 3476 194652 3528
rect 195612 3476 195664 3528
rect 198648 3476 198700 3528
rect 199108 3476 199160 3528
rect 202788 3476 202840 3528
rect 203892 3476 203944 3528
rect 205548 3476 205600 3528
rect 206192 3476 206244 3528
rect 206928 3476 206980 3528
rect 207388 3476 207440 3528
rect 211068 3476 211120 3528
rect 212172 3476 212224 3528
rect 215208 3476 215260 3528
rect 216864 3476 216916 3528
rect 217968 3476 218020 3528
rect 219256 3476 219308 3528
rect 220084 3476 220136 3528
rect 221556 3476 221608 3528
rect 222844 3476 222896 3528
rect 223948 3476 224000 3528
rect 227628 3476 227680 3528
rect 229836 3476 229888 3528
rect 233148 3476 233200 3528
rect 235816 3476 235868 3528
rect 240784 3476 240836 3528
rect 244096 3476 244148 3528
rect 246948 3476 247000 3528
rect 251180 3476 251232 3528
rect 256608 3476 256660 3528
rect 261760 3476 261812 3528
rect 269028 3476 269080 3528
rect 274824 3476 274876 3528
rect 289728 3476 289780 3528
rect 297272 3476 297324 3528
rect 299296 3476 299348 3528
rect 306748 3476 306800 3528
rect 307668 3476 307720 3528
rect 316224 3476 316276 3528
rect 321468 3476 321520 3528
rect 331588 3476 331640 3528
rect 335268 3612 335320 3664
rect 345756 3612 345808 3664
rect 346216 3612 346268 3664
rect 358728 3612 358780 3664
rect 361488 3748 361540 3800
rect 374092 3748 374144 3800
rect 380808 3748 380860 3800
rect 395344 3748 395396 3800
rect 395988 3748 396040 3800
rect 411904 3748 411956 3800
rect 415308 3748 415360 3800
rect 432052 3748 432104 3800
rect 437296 3748 437348 3800
rect 455696 3748 455748 3800
rect 460848 3748 460900 3800
rect 481732 3748 481784 3800
rect 484216 3748 484268 3800
rect 506480 3748 506532 3800
rect 513288 3748 513340 3800
rect 538404 3748 538456 3800
rect 545028 3748 545080 3800
rect 572720 3748 572772 3800
rect 362776 3680 362828 3732
rect 376484 3680 376536 3732
rect 376668 3680 376720 3732
rect 390652 3680 390704 3732
rect 391848 3680 391900 3732
rect 407212 3680 407264 3732
rect 411168 3680 411220 3732
rect 428464 3680 428516 3732
rect 431776 3680 431828 3732
rect 450912 3680 450964 3732
rect 452476 3680 452528 3732
rect 453948 3680 454000 3732
rect 474556 3680 474608 3732
rect 474648 3680 474700 3732
rect 495900 3680 495952 3732
rect 496728 3680 496780 3732
rect 520740 3680 520792 3732
rect 526996 3680 527048 3732
rect 552664 3680 552716 3732
rect 553308 3680 553360 3732
rect 582196 3680 582248 3732
rect 371700 3612 371752 3664
rect 375288 3612 375340 3664
rect 389456 3612 389508 3664
rect 390468 3612 390520 3664
rect 406016 3612 406068 3664
rect 407028 3612 407080 3664
rect 423772 3612 423824 3664
rect 427728 3612 427780 3664
rect 446220 3612 446272 3664
rect 448336 3612 448388 3664
rect 468668 3612 468720 3664
rect 474464 3612 474516 3664
rect 497096 3612 497148 3664
rect 498108 3612 498160 3664
rect 521844 3612 521896 3664
rect 522948 3612 523000 3664
rect 549076 3612 549128 3664
rect 550548 3612 550600 3664
rect 578608 3612 578660 3664
rect 338028 3544 338080 3596
rect 349252 3544 349304 3596
rect 353208 3544 353260 3596
rect 365812 3544 365864 3596
rect 368296 3544 368348 3596
rect 381176 3544 381228 3596
rect 383568 3544 383620 3596
rect 398932 3544 398984 3596
rect 400036 3544 400088 3596
rect 415492 3544 415544 3596
rect 420828 3544 420880 3596
rect 439136 3544 439188 3596
rect 442816 3544 442868 3596
rect 462780 3544 462832 3596
rect 464988 3544 465040 3596
rect 486424 3544 486476 3596
rect 489828 3544 489880 3596
rect 513564 3544 513616 3596
rect 520188 3544 520240 3596
rect 545488 3544 545540 3596
rect 549168 3544 549220 3596
rect 577412 3544 577464 3596
rect 342168 3476 342220 3528
rect 344928 3476 344980 3528
rect 356336 3476 356388 3528
rect 361120 3476 361172 3528
rect 73804 3408 73856 3460
rect 74448 3408 74500 3460
rect 131764 3408 131816 3460
rect 132408 3408 132460 3460
rect 135260 3408 135312 3460
rect 136548 3408 136600 3460
rect 155408 3408 155460 3460
rect 155868 3408 155920 3460
rect 195980 3408 196032 3460
rect 196808 3408 196860 3460
rect 216588 3408 216640 3460
rect 218060 3408 218112 3460
rect 224868 3408 224920 3460
rect 227536 3408 227588 3460
rect 231768 3408 231820 3460
rect 234620 3408 234672 3460
rect 241428 3408 241480 3460
rect 245200 3408 245252 3460
rect 249708 3408 249760 3460
rect 253480 3408 253532 3460
rect 259368 3408 259420 3460
rect 264152 3408 264204 3460
rect 267556 3408 267608 3460
rect 273628 3408 273680 3460
rect 277216 3408 277268 3460
rect 284300 3408 284352 3460
rect 296628 3408 296680 3460
rect 304356 3408 304408 3460
rect 304816 3408 304868 3460
rect 313832 3408 313884 3460
rect 314476 3408 314528 3460
rect 324412 3408 324464 3460
rect 325700 3408 325752 3460
rect 336280 3408 336332 3460
rect 336556 3408 336608 3460
rect 348056 3408 348108 3460
rect 351828 3408 351880 3460
rect 300676 3340 300728 3392
rect 309048 3340 309100 3392
rect 319996 3340 320048 3392
rect 330392 3340 330444 3392
rect 333796 3340 333848 3392
rect 344560 3340 344612 3392
rect 357256 3340 357308 3392
rect 370596 3476 370648 3528
rect 379336 3476 379388 3528
rect 394240 3476 394292 3528
rect 397368 3476 397420 3528
rect 413100 3476 413152 3528
rect 415216 3476 415268 3528
rect 433248 3476 433300 3528
rect 437388 3476 437440 3528
rect 456892 3476 456944 3528
rect 458088 3476 458140 3528
rect 479340 3476 479392 3528
rect 480168 3476 480220 3528
rect 502984 3476 503036 3528
rect 506388 3476 506440 3528
rect 531320 3476 531372 3528
rect 543556 3476 543608 3528
rect 571524 3476 571576 3528
rect 364616 3408 364668 3460
rect 368388 3408 368440 3460
rect 382372 3408 382424 3460
rect 388996 3408 389048 3460
rect 404820 3408 404872 3460
rect 405556 3408 405608 3460
rect 422576 3408 422628 3460
rect 426256 3408 426308 3460
rect 445024 3408 445076 3460
rect 449900 3408 449952 3460
rect 80888 3272 80940 3324
rect 81348 3272 81400 3324
rect 85672 3272 85724 3324
rect 86776 3272 86828 3324
rect 89168 3272 89220 3324
rect 89628 3272 89680 3324
rect 126980 3272 127032 3324
rect 130384 3272 130436 3324
rect 220728 3272 220780 3324
rect 222752 3272 222804 3324
rect 252468 3272 252520 3324
rect 257068 3272 257120 3324
rect 260748 3272 260800 3324
rect 265348 3272 265400 3324
rect 271788 3272 271840 3324
rect 277124 3272 277176 3324
rect 278688 3272 278740 3324
rect 285404 3272 285456 3324
rect 288256 3272 288308 3324
rect 296076 3272 296128 3324
rect 298008 3272 298060 3324
rect 305552 3272 305604 3324
rect 350356 3272 350408 3324
rect 362316 3272 362368 3324
rect 84476 3204 84528 3256
rect 85488 3204 85540 3256
rect 208308 3204 208360 3256
rect 209780 3204 209832 3256
rect 245568 3204 245620 3256
rect 230388 3136 230440 3188
rect 233424 3136 233476 3188
rect 234528 3136 234580 3188
rect 237012 3136 237064 3188
rect 240048 3136 240100 3188
rect 242900 3136 242952 3188
rect 246304 3136 246356 3188
rect 247592 3136 247644 3188
rect 250996 3204 251048 3256
rect 254676 3204 254728 3256
rect 340788 3204 340840 3256
rect 351644 3204 351696 3256
rect 357348 3204 357400 3256
rect 369400 3340 369452 3392
rect 372528 3340 372580 3392
rect 385960 3340 386012 3392
rect 386328 3340 386380 3392
rect 401324 3340 401376 3392
rect 364248 3272 364300 3324
rect 377680 3272 377732 3324
rect 389088 3272 389140 3324
rect 403624 3272 403676 3324
rect 362868 3204 362920 3256
rect 375288 3204 375340 3256
rect 379428 3204 379480 3256
rect 393044 3204 393096 3256
rect 401508 3204 401560 3256
rect 405648 3272 405700 3324
rect 248788 3136 248840 3188
rect 264244 3136 264296 3188
rect 266544 3136 266596 3188
rect 273168 3136 273220 3188
rect 279516 3136 279568 3188
rect 369768 3136 369820 3188
rect 383568 3136 383620 3188
rect 387708 3136 387760 3188
rect 402520 3136 402572 3188
rect 408316 3136 408368 3188
rect 413928 3340 413980 3392
rect 430856 3340 430908 3392
rect 445668 3340 445720 3392
rect 409788 3272 409840 3324
rect 426164 3272 426216 3324
rect 431868 3272 431920 3324
rect 449716 3272 449768 3324
rect 473452 3408 473504 3460
rect 491208 3408 491260 3460
rect 514760 3408 514812 3460
rect 517336 3408 517388 3460
rect 543188 3408 543240 3460
rect 551928 3408 551980 3460
rect 581000 3408 581052 3460
rect 465172 3340 465224 3392
rect 469128 3340 469180 3392
rect 489920 3340 489972 3392
rect 500868 3340 500920 3392
rect 525432 3340 525484 3392
rect 527088 3340 527140 3392
rect 553768 3340 553820 3392
rect 469864 3272 469916 3324
rect 471888 3272 471940 3324
rect 493508 3272 493560 3324
rect 503628 3272 503680 3324
rect 527824 3272 527876 3324
rect 532608 3272 532660 3324
rect 559748 3272 559800 3324
rect 417884 3204 417936 3256
rect 418068 3204 418120 3256
rect 435548 3204 435600 3256
rect 440148 3204 440200 3256
rect 459192 3204 459244 3256
rect 462228 3204 462280 3256
rect 482836 3204 482888 3256
rect 488448 3204 488500 3256
rect 511264 3204 511316 3256
rect 511908 3204 511960 3256
rect 536104 3204 536156 3256
rect 536748 3204 536800 3256
rect 563244 3204 563296 3256
rect 378048 3068 378100 3120
rect 391848 3068 391900 3120
rect 393228 3068 393280 3120
rect 408408 3068 408460 3120
rect 421380 3136 421432 3188
rect 424876 3136 424928 3188
rect 424968 3068 425020 3120
rect 433156 3136 433208 3188
rect 452108 3136 452160 3188
rect 452568 3136 452620 3188
rect 455328 3136 455380 3188
rect 475752 3136 475804 3188
rect 478788 3136 478840 3188
rect 500592 3136 500644 3188
rect 517428 3136 517480 3188
rect 541992 3136 542044 3188
rect 547788 3136 547840 3188
rect 575112 3136 575164 3188
rect 442632 3068 442684 3120
rect 448428 3068 448480 3120
rect 467472 3068 467524 3120
rect 467748 3068 467800 3120
rect 488816 3068 488868 3120
rect 500776 3068 500828 3120
rect 524236 3068 524288 3120
rect 540888 3068 540940 3120
rect 568028 3068 568080 3120
rect 143540 3000 143592 3052
rect 144644 3000 144696 3052
rect 150624 3000 150676 3052
rect 151728 3000 151780 3052
rect 263508 3000 263560 3052
rect 268844 3000 268896 3052
rect 291108 3000 291160 3052
rect 298468 3000 298520 3052
rect 402888 3000 402940 3052
rect 418988 3000 419040 3052
rect 419448 3000 419500 3052
rect 436744 3000 436796 3052
rect 438768 3000 438820 3052
rect 458088 3000 458140 3052
rect 495348 3000 495400 3052
rect 518348 3000 518400 3052
rect 538128 3000 538180 3052
rect 564440 3000 564492 3052
rect 583392 3000 583444 3052
rect 25320 2932 25372 2984
rect 26148 2932 26200 2984
rect 83280 2932 83332 2984
rect 84108 2932 84160 2984
rect 213828 2932 213880 2984
rect 215668 2932 215720 2984
rect 224776 2932 224828 2984
rect 226340 2932 226392 2984
rect 270408 2932 270460 2984
rect 276020 2932 276072 2984
rect 280068 2932 280120 2984
rect 286600 2932 286652 2984
rect 404268 2932 404320 2984
rect 420184 2932 420236 2984
rect 423588 2932 423640 2984
rect 441528 2932 441580 2984
rect 442908 2932 442960 2984
rect 255228 2864 255280 2916
rect 259460 2864 259512 2916
rect 288348 2864 288400 2916
rect 294880 2864 294932 2916
rect 426348 2864 426400 2916
rect 443828 2864 443880 2916
rect 447048 2932 447100 2984
rect 466276 2932 466328 2984
rect 533988 2932 534040 2984
rect 560852 2932 560904 2984
rect 461584 2864 461636 2916
rect 531228 2864 531280 2916
rect 557356 2864 557408 2916
rect 436008 2796 436060 2848
rect 454500 2796 454552 2848
rect 472256 2796 472308 2848
rect 524328 2796 524380 2848
rect 550272 2796 550324 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700534 40540 703520
rect 72988 700670 73016 703520
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 40500 700528 40552 700534
rect 40500 700470 40552 700476
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 105464 699718 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 170324 700466 170352 703520
rect 170312 700460 170364 700466
rect 170312 700402 170364 700408
rect 180064 700460 180116 700466
rect 180064 700402 180116 700408
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 106200 674218 106228 699654
rect 180076 674354 180104 700402
rect 202800 700126 202828 703520
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 218992 700058 219020 703520
rect 233148 700596 233200 700602
rect 233148 700538 233200 700544
rect 218980 700052 219032 700058
rect 218980 699994 219032 700000
rect 219348 696992 219400 696998
rect 219348 696934 219400 696940
rect 180064 674348 180116 674354
rect 180064 674290 180116 674296
rect 106188 674212 106240 674218
rect 106188 674154 106240 674160
rect 219360 673470 219388 696934
rect 223488 683188 223540 683194
rect 223488 683130 223540 683136
rect 218152 673464 218204 673470
rect 218152 673406 218204 673412
rect 219348 673464 219400 673470
rect 223500 673454 223528 683130
rect 227536 674144 227588 674150
rect 227536 674086 227588 674092
rect 219348 673406 219400 673412
rect 223224 673426 223528 673454
rect 204352 673396 204404 673402
rect 204352 673338 204404 673344
rect 67916 673328 67968 673334
rect 67916 673270 67968 673276
rect 5172 673192 5224 673198
rect 5172 673134 5224 673140
rect 5080 673124 5132 673130
rect 5080 673066 5132 673072
rect 4988 672920 5040 672926
rect 4988 672862 5040 672868
rect 4804 672172 4856 672178
rect 4804 672114 4856 672120
rect 3056 672036 3108 672042
rect 3056 671978 3108 671984
rect 3068 671265 3096 671978
rect 3054 671256 3110 671265
rect 3054 671191 3110 671200
rect 3884 670472 3936 670478
rect 3884 670414 3936 670420
rect 3792 668704 3844 668710
rect 3792 668646 3844 668652
rect 3424 668636 3476 668642
rect 3424 668578 3476 668584
rect 3240 658232 3292 658238
rect 3238 658200 3240 658209
rect 3292 658200 3294 658209
rect 3238 658135 3294 658144
rect 3332 632188 3384 632194
rect 3332 632130 3384 632136
rect 3344 632097 3372 632130
rect 3330 632088 3386 632097
rect 3330 632023 3386 632032
rect 2964 619336 3016 619342
rect 2964 619278 3016 619284
rect 2976 619177 3004 619278
rect 2962 619168 3018 619177
rect 2962 619103 3018 619112
rect 2872 607164 2924 607170
rect 2872 607106 2924 607112
rect 2884 606121 2912 607106
rect 2870 606112 2926 606121
rect 2870 606047 2926 606056
rect 3148 580508 3200 580514
rect 3148 580450 3200 580456
rect 3160 580009 3188 580450
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 3332 554736 3384 554742
rect 3332 554678 3384 554684
rect 3344 553897 3372 554678
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3240 528556 3292 528562
rect 3240 528498 3292 528504
rect 3252 527921 3280 528498
rect 3238 527912 3294 527921
rect 3238 527847 3294 527856
rect 2780 515636 2832 515642
rect 2780 515578 2832 515584
rect 2792 514865 2820 515578
rect 2778 514856 2834 514865
rect 2778 514791 2834 514800
rect 3332 502308 3384 502314
rect 3332 502250 3384 502256
rect 3344 501809 3372 502250
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3332 476060 3384 476066
rect 3332 476002 3384 476008
rect 3344 475697 3372 476002
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 2780 463480 2832 463486
rect 2780 463422 2832 463428
rect 2792 462641 2820 463422
rect 2778 462632 2834 462641
rect 2778 462567 2834 462576
rect 2964 449608 3016 449614
rect 2962 449576 2964 449585
rect 3016 449576 3018 449585
rect 2962 449511 3018 449520
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3332 371612 3384 371618
rect 3332 371554 3384 371560
rect 3344 371385 3372 371554
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 2832 358456 2834 358465
rect 2778 358391 2834 358400
rect 2964 346384 3016 346390
rect 2964 346326 3016 346332
rect 2976 345409 3004 346326
rect 2962 345400 3018 345409
rect 2962 345335 3018 345344
rect 3240 320068 3292 320074
rect 3240 320010 3292 320016
rect 3252 319297 3280 320010
rect 3238 319288 3294 319297
rect 3238 319223 3294 319232
rect 3332 306264 3384 306270
rect 3330 306232 3332 306241
rect 3384 306232 3386 306241
rect 3330 306167 3386 306176
rect 3240 267708 3292 267714
rect 3240 267650 3292 267656
rect 3252 267209 3280 267650
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3332 255264 3384 255270
rect 3332 255206 3384 255212
rect 3344 254153 3372 255206
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 2780 241120 2832 241126
rect 2778 241088 2780 241097
rect 2832 241088 2834 241097
rect 2778 241023 2834 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3332 202836 3384 202842
rect 3332 202778 3384 202784
rect 3344 201929 3372 202778
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 2780 136876 2832 136882
rect 2780 136818 2832 136824
rect 2792 136785 2820 136818
rect 2778 136776 2834 136785
rect 2778 136711 2834 136720
rect 2964 111172 3016 111178
rect 2964 111114 3016 111120
rect 2976 110673 3004 111114
rect 2962 110664 3018 110673
rect 2962 110599 3018 110608
rect 3240 97980 3292 97986
rect 3240 97922 3292 97928
rect 3252 97617 3280 97922
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2688 47796 2740 47802
rect 2688 47738 2740 47744
rect 1308 47592 1360 47598
rect 1308 47534 1360 47540
rect 1320 3534 1348 47534
rect 2700 3534 2728 47738
rect 2780 32972 2832 32978
rect 2780 32914 2832 32920
rect 2792 32473 2820 32914
rect 2778 32464 2834 32473
rect 2778 32399 2834 32408
rect 3436 6497 3464 668578
rect 3700 668432 3752 668438
rect 3700 668374 3752 668380
rect 3608 668296 3660 668302
rect 3608 668238 3660 668244
rect 3516 668228 3568 668234
rect 3516 668170 3568 668176
rect 3528 84697 3556 668170
rect 3620 188873 3648 668238
rect 3712 293185 3740 668374
rect 3804 397497 3832 668646
rect 3896 566953 3924 670414
rect 3882 566944 3938 566953
rect 3882 566879 3938 566888
rect 3790 397488 3846 397497
rect 3790 397423 3846 397432
rect 3698 293176 3754 293185
rect 3698 293111 3754 293120
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3608 150408 3660 150414
rect 3608 150350 3660 150356
rect 3620 149841 3648 150350
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 4816 136882 4844 672114
rect 4896 668364 4948 668370
rect 4896 668306 4948 668312
rect 4908 241126 4936 668306
rect 5000 358494 5028 672862
rect 5092 463486 5120 673066
rect 5184 515642 5212 673134
rect 7840 672716 7892 672722
rect 7840 672658 7892 672664
rect 7748 672104 7800 672110
rect 7748 672046 7800 672052
rect 7656 670880 7708 670886
rect 6182 670848 6238 670857
rect 7656 670822 7708 670828
rect 6182 670783 6238 670792
rect 5172 515636 5224 515642
rect 5172 515578 5224 515584
rect 5080 463480 5132 463486
rect 5080 463422 5132 463428
rect 4988 358488 5040 358494
rect 4988 358430 5040 358436
rect 4896 241120 4948 241126
rect 4896 241062 4948 241068
rect 4804 136876 4856 136882
rect 4804 136818 4856 136824
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71664 3568 71670
rect 3514 71632 3516 71641
rect 3568 71632 3570 71641
rect 3514 71567 3570 71576
rect 4068 48204 4120 48210
rect 4068 48146 4120 48152
rect 3976 47660 4028 47666
rect 3976 47602 4028 47608
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3528 19417 3556 20606
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3988 16574 4016 47602
rect 3896 16546 4016 16574
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 584 480 612 3470
rect 1688 480 1716 3470
rect 2884 480 2912 3538
rect 3896 3482 3924 16546
rect 4080 6914 4108 48146
rect 5448 47864 5500 47870
rect 5448 47806 5500 47812
rect 5460 6914 5488 47806
rect 6196 32978 6224 670783
rect 6368 670676 6420 670682
rect 6368 670618 6420 670624
rect 6276 668772 6328 668778
rect 6276 668714 6328 668720
rect 6288 449614 6316 668714
rect 6380 658238 6408 670618
rect 7564 668024 7616 668030
rect 7564 667966 7616 667972
rect 6368 658232 6420 658238
rect 6368 658174 6420 658180
rect 6276 449608 6328 449614
rect 6276 449550 6328 449556
rect 6828 47932 6880 47938
rect 6828 47874 6880 47880
rect 6184 32972 6236 32978
rect 6184 32914 6236 32920
rect 6840 6914 6868 47874
rect 7576 45558 7604 667966
rect 7668 111178 7696 670822
rect 7760 150414 7788 672046
rect 7852 306270 7880 672658
rect 11888 672648 11940 672654
rect 11888 672590 11940 672596
rect 11702 672480 11758 672489
rect 11702 672415 11758 672424
rect 10322 672208 10378 672217
rect 10322 672143 10378 672152
rect 7932 671356 7984 671362
rect 7932 671298 7984 671304
rect 7944 371618 7972 671298
rect 9036 671288 9088 671294
rect 9036 671230 9088 671236
rect 8942 670984 8998 670993
rect 8942 670919 8998 670928
rect 8024 670608 8076 670614
rect 8024 670550 8076 670556
rect 8036 632194 8064 670550
rect 8024 632188 8076 632194
rect 8024 632130 8076 632136
rect 7932 371612 7984 371618
rect 7932 371554 7984 371560
rect 7840 306264 7892 306270
rect 7840 306206 7892 306212
rect 7748 150408 7800 150414
rect 7748 150350 7800 150356
rect 7656 111172 7708 111178
rect 7656 111114 7708 111120
rect 8956 71670 8984 670919
rect 9048 320074 9076 671230
rect 9220 670404 9272 670410
rect 9220 670346 9272 670352
rect 9128 670336 9180 670342
rect 9128 670278 9180 670284
rect 9140 580514 9168 670278
rect 9232 619342 9260 670346
rect 9220 619336 9272 619342
rect 9220 619278 9272 619284
rect 9128 580508 9180 580514
rect 9128 580450 9180 580456
rect 9036 320068 9088 320074
rect 9036 320010 9088 320016
rect 8944 71664 8996 71670
rect 8944 71606 8996 71612
rect 8208 48136 8260 48142
rect 8208 48078 8260 48084
rect 7564 45552 7616 45558
rect 7564 45494 7616 45500
rect 3988 6886 4108 6914
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 3988 3602 4016 6886
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3896 3454 4108 3482
rect 4080 480 4108 3454
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 8220 3534 8248 48078
rect 9588 47728 9640 47734
rect 9588 47670 9640 47676
rect 9600 3534 9628 47670
rect 10336 20670 10364 672143
rect 10692 671968 10744 671974
rect 10692 671910 10744 671916
rect 10416 671152 10468 671158
rect 10416 671094 10468 671100
rect 10428 267714 10456 671094
rect 10600 670064 10652 670070
rect 10600 670006 10652 670012
rect 10508 668568 10560 668574
rect 10508 668510 10560 668516
rect 10520 346390 10548 668510
rect 10612 528562 10640 670006
rect 10704 607170 10732 671910
rect 10692 607164 10744 607170
rect 10692 607106 10744 607112
rect 10600 528556 10652 528562
rect 10600 528498 10652 528504
rect 10508 346384 10560 346390
rect 10508 346326 10560 346332
rect 10416 267708 10468 267714
rect 10416 267650 10468 267656
rect 11716 97986 11744 672415
rect 11796 671084 11848 671090
rect 11796 671026 11848 671032
rect 11808 215286 11836 671026
rect 11900 255270 11928 672590
rect 13268 672512 13320 672518
rect 13268 672454 13320 672460
rect 13082 672344 13138 672353
rect 13082 672279 13138 672288
rect 12072 671560 12124 671566
rect 12072 671502 12124 671508
rect 11980 669860 12032 669866
rect 11980 669802 12032 669808
rect 11992 411262 12020 669802
rect 12084 476066 12112 671502
rect 12164 670268 12216 670274
rect 12164 670210 12216 670216
rect 12176 554742 12204 670210
rect 12164 554736 12216 554742
rect 12164 554678 12216 554684
rect 12072 476060 12124 476066
rect 12072 476002 12124 476008
rect 11980 411256 12032 411262
rect 11980 411198 12032 411204
rect 11888 255264 11940 255270
rect 11888 255206 11940 255212
rect 11796 215280 11848 215286
rect 11796 215222 11848 215228
rect 11704 97980 11756 97986
rect 11704 97922 11756 97928
rect 13096 59362 13124 672279
rect 13176 670948 13228 670954
rect 13176 670890 13228 670896
rect 13188 164218 13216 670890
rect 13280 202842 13308 672454
rect 13452 671696 13504 671702
rect 13452 671638 13504 671644
rect 13360 671492 13412 671498
rect 13360 671434 13412 671440
rect 13372 423638 13400 671434
rect 13464 502314 13492 671638
rect 58532 670812 58584 670818
rect 58532 670754 58584 670760
rect 44456 670744 44508 670750
rect 35070 670712 35126 670721
rect 44456 670686 44508 670692
rect 35070 670647 35126 670656
rect 35084 669868 35112 670647
rect 44468 669868 44496 670686
rect 58544 669868 58572 670754
rect 67928 669868 67956 673270
rect 180616 673260 180668 673266
rect 180616 673202 180668 673208
rect 147772 673056 147824 673062
rect 147772 672998 147824 673004
rect 138388 672988 138440 672994
rect 138388 672930 138440 672936
rect 124312 672852 124364 672858
rect 124312 672794 124364 672800
rect 119528 672784 119580 672790
rect 119528 672726 119580 672732
rect 105452 672580 105504 672586
rect 105452 672522 105504 672528
rect 81992 672444 82044 672450
rect 81992 672386 82044 672392
rect 77300 672240 77352 672246
rect 77300 672182 77352 672188
rect 77312 669868 77340 672182
rect 82004 669868 82032 672386
rect 91376 672376 91428 672382
rect 91376 672318 91428 672324
rect 86684 671016 86736 671022
rect 86684 670958 86736 670964
rect 86696 669868 86724 670958
rect 91388 669868 91416 672318
rect 96068 672308 96120 672314
rect 96068 672250 96120 672256
rect 96080 669868 96108 672250
rect 105464 669868 105492 672522
rect 114836 671220 114888 671226
rect 114836 671162 114888 671168
rect 114848 669868 114876 671162
rect 119540 669868 119568 672726
rect 124324 669868 124352 672794
rect 138400 669868 138428 672930
rect 143080 671424 143132 671430
rect 143080 671366 143132 671372
rect 143092 669868 143120 671366
rect 147784 669868 147812 672998
rect 161848 671628 161900 671634
rect 161848 671570 161900 671576
rect 157064 669928 157116 669934
rect 157116 669876 157182 669882
rect 157064 669870 157182 669876
rect 157076 669854 157182 669870
rect 161860 669868 161888 671570
rect 175924 670132 175976 670138
rect 175924 670074 175976 670080
rect 166816 669996 166868 670002
rect 166816 669938 166868 669944
rect 171600 669996 171652 670002
rect 171600 669938 171652 669944
rect 166828 669882 166856 669938
rect 171612 669882 171640 669938
rect 166566 669854 166856 669882
rect 171258 669854 171640 669882
rect 175936 669868 175964 670074
rect 180628 669868 180656 673202
rect 199384 671900 199436 671906
rect 199384 671842 199436 671848
rect 190000 671764 190052 671770
rect 190000 671706 190052 671712
rect 185308 670200 185360 670206
rect 185308 670142 185360 670148
rect 185320 669868 185348 670142
rect 190012 669868 190040 671706
rect 199396 669868 199424 671842
rect 204076 670540 204128 670546
rect 204076 670482 204128 670488
rect 204088 669868 204116 670482
rect 204364 670478 204392 673338
rect 213460 671832 213512 671838
rect 213460 671774 213512 671780
rect 204352 670472 204404 670478
rect 204352 670414 204404 670420
rect 208768 670472 208820 670478
rect 208768 670414 208820 670420
rect 208780 669868 208808 670414
rect 213472 669868 213500 671774
rect 218164 669868 218192 673406
rect 223224 669882 223252 673426
rect 222870 669854 223252 669882
rect 227548 669868 227576 674086
rect 233160 673470 233188 700538
rect 235184 699854 235212 703520
rect 246948 700868 247000 700874
rect 246948 700810 247000 700816
rect 237288 700460 237340 700466
rect 237288 700402 237340 700408
rect 235172 699848 235224 699854
rect 235172 699790 235224 699796
rect 232320 673464 232372 673470
rect 232320 673406 232372 673412
rect 233148 673464 233200 673470
rect 233148 673406 233200 673412
rect 232332 669868 232360 673406
rect 237300 669882 237328 700402
rect 238024 699848 238076 699854
rect 238024 699790 238076 699796
rect 238036 674490 238064 699790
rect 238024 674484 238076 674490
rect 238024 674426 238076 674432
rect 241704 674280 241756 674286
rect 241704 674222 241756 674228
rect 237038 669854 237328 669882
rect 241716 669868 241744 674222
rect 246960 673454 246988 700810
rect 251088 700800 251140 700806
rect 251088 700742 251140 700748
rect 246776 673426 246988 673454
rect 246776 669882 246804 673426
rect 246422 669854 246804 669882
rect 251100 669868 251128 700742
rect 266268 700256 266320 700262
rect 266268 700198 266320 700204
rect 260748 700188 260800 700194
rect 260748 700130 260800 700136
rect 256608 676864 256660 676870
rect 256608 676806 256660 676812
rect 256620 673470 256648 676806
rect 255780 673464 255832 673470
rect 255780 673406 255832 673412
rect 256608 673464 256660 673470
rect 256608 673406 256660 673412
rect 255792 669868 255820 673406
rect 260760 669882 260788 700130
rect 266280 673470 266308 700198
rect 267660 699854 267688 703520
rect 280068 699984 280120 699990
rect 280068 699926 280120 699932
rect 274548 699916 274600 699922
rect 274548 699858 274600 699864
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 269856 674416 269908 674422
rect 269856 674358 269908 674364
rect 265164 673464 265216 673470
rect 265164 673406 265216 673412
rect 266268 673464 266320 673470
rect 266268 673406 266320 673412
rect 260498 669854 260788 669882
rect 265176 669868 265204 673406
rect 269868 669868 269896 674358
rect 274560 669868 274588 699858
rect 280080 673470 280108 699926
rect 283852 699786 283880 703520
rect 288440 699848 288492 699854
rect 288440 699790 288492 699796
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 283932 674552 283984 674558
rect 283932 674494 283984 674500
rect 279240 673464 279292 673470
rect 279240 673406 279292 673412
rect 280068 673464 280120 673470
rect 280068 673406 280120 673412
rect 279252 669868 279280 673406
rect 283944 669868 283972 674494
rect 288452 669882 288480 699790
rect 292580 699780 292632 699786
rect 292580 699722 292632 699728
rect 292592 692774 292620 699722
rect 292592 692746 292896 692774
rect 292868 669882 292896 692746
rect 299492 674558 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 320180 701004 320232 701010
rect 320180 700946 320232 700952
rect 316040 700936 316092 700942
rect 316040 700878 316092 700884
rect 302240 700120 302292 700126
rect 302240 700062 302292 700068
rect 299480 674552 299532 674558
rect 299480 674494 299532 674500
rect 298008 674484 298060 674490
rect 298008 674426 298060 674432
rect 288452 669854 288650 669882
rect 292868 669854 293342 669882
rect 298020 669868 298048 674426
rect 302252 669882 302280 700062
rect 306380 700052 306432 700058
rect 306380 699994 306432 700000
rect 306392 692774 306420 699994
rect 316052 692774 316080 700878
rect 320192 692774 320220 700946
rect 329840 700664 329892 700670
rect 329840 700606 329892 700612
rect 331864 700664 331916 700670
rect 331864 700606 331916 700612
rect 329852 692774 329880 700606
rect 306392 692746 307064 692774
rect 316052 692746 316448 692774
rect 320192 692746 321048 692774
rect 329852 692746 330432 692774
rect 307036 669882 307064 692746
rect 312084 674348 312136 674354
rect 312084 674290 312136 674296
rect 302252 669854 302726 669882
rect 307036 669854 307418 669882
rect 312096 669868 312124 674290
rect 316420 669882 316448 692746
rect 321020 669882 321048 692746
rect 326160 674212 326212 674218
rect 326160 674154 326212 674160
rect 316420 669854 316802 669882
rect 321020 669854 321494 669882
rect 326172 669868 326200 674154
rect 330404 669882 330432 692746
rect 331876 676870 331904 700606
rect 332520 699922 332548 703520
rect 335360 700732 335412 700738
rect 335360 700674 335412 700680
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 331864 676864 331916 676870
rect 331864 676806 331916 676812
rect 335372 669882 335400 700674
rect 339500 700528 339552 700534
rect 339500 700470 339552 700476
rect 339512 692774 339540 700470
rect 345020 700324 345072 700330
rect 345020 700266 345072 700272
rect 339512 692746 340000 692774
rect 339972 669882 340000 692746
rect 330404 669854 330878 669882
rect 335372 669854 335570 669882
rect 339972 669854 340354 669882
rect 345032 669868 345060 700266
rect 348804 699990 348832 703520
rect 349160 700392 349212 700398
rect 349160 700334 349212 700340
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 349172 692774 349200 700334
rect 364996 699718 365024 703520
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 429856 700670 429884 703520
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 429844 700664 429896 700670
rect 429844 700606 429896 700612
rect 494808 700330 494836 703520
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 443644 700324 443696 700330
rect 443644 700266 443696 700272
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 363604 699712 363656 699718
rect 363604 699654 363656 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 349172 692746 349384 692774
rect 349356 669882 349384 692746
rect 353944 683256 353996 683262
rect 353944 683198 353996 683204
rect 353956 669882 353984 683198
rect 363616 674422 363644 699654
rect 363604 674416 363656 674422
rect 363604 674358 363656 674364
rect 443656 674286 443684 700266
rect 559668 699718 559696 703520
rect 555424 699712 555476 699718
rect 555424 699654 555476 699660
rect 559656 699712 559708 699718
rect 559656 699654 559708 699660
rect 443644 674280 443696 674286
rect 443644 674222 443696 674228
rect 555436 674150 555464 699654
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 555424 674144 555476 674150
rect 555424 674086 555476 674092
rect 391940 673396 391992 673402
rect 391940 673338 391992 673344
rect 359464 673328 359516 673334
rect 359464 673270 359516 673276
rect 359476 670682 359504 673270
rect 363788 672036 363840 672042
rect 363788 671978 363840 671984
rect 359096 670676 359148 670682
rect 359096 670618 359148 670624
rect 359464 670676 359516 670682
rect 359464 670618 359516 670624
rect 349356 669854 349738 669882
rect 353956 669854 354430 669882
rect 359108 669868 359136 670618
rect 363800 669868 363828 671978
rect 373172 671968 373224 671974
rect 373172 671910 373224 671916
rect 368480 670608 368532 670614
rect 368480 670550 368532 670556
rect 368492 669868 368520 670550
rect 373184 669868 373212 671910
rect 377864 670404 377916 670410
rect 377864 670346 377916 670352
rect 377876 669868 377904 670346
rect 382556 670336 382608 670342
rect 382556 670278 382608 670284
rect 382568 669868 382596 670278
rect 387248 670268 387300 670274
rect 387248 670210 387300 670216
rect 387260 669868 387288 670210
rect 391952 669868 391980 673338
rect 555516 673260 555568 673266
rect 555516 673202 555568 673208
rect 406016 673192 406068 673198
rect 406016 673134 406068 673140
rect 401324 671696 401376 671702
rect 401324 671638 401376 671644
rect 396356 670064 396408 670070
rect 396356 670006 396408 670012
rect 396368 669882 396396 670006
rect 396368 669854 396658 669882
rect 401336 669868 401364 671638
rect 406028 669868 406056 673134
rect 420092 673124 420144 673130
rect 420092 673066 420144 673072
rect 410708 671560 410760 671566
rect 410708 671502 410760 671508
rect 410720 669868 410748 671502
rect 415308 670064 415360 670070
rect 415308 670006 415360 670012
rect 415320 669882 415348 670006
rect 415320 669854 415426 669882
rect 420104 669868 420132 673066
rect 448336 672920 448388 672926
rect 448336 672862 448388 672868
rect 424784 671492 424836 671498
rect 424784 671434 424836 671440
rect 424796 669868 424824 671434
rect 438860 671356 438912 671362
rect 438860 671298 438912 671304
rect 433892 670064 433944 670070
rect 433892 670006 433944 670012
rect 433904 669882 433932 670006
rect 429212 669866 429502 669882
rect 429200 669860 429502 669866
rect 429252 669854 429502 669860
rect 433904 669854 434194 669882
rect 438872 669868 438900 671298
rect 443288 669866 443578 669882
rect 448348 669868 448376 672862
rect 462412 672716 462464 672722
rect 462412 672658 462464 672664
rect 453028 671288 453080 671294
rect 453028 671230 453080 671236
rect 453040 669868 453068 671230
rect 457456 669866 457746 669882
rect 462424 669868 462452 672658
rect 476488 672648 476540 672654
rect 476488 672590 476540 672596
rect 467104 671152 467156 671158
rect 467104 671094 467156 671100
rect 467116 669868 467144 671094
rect 471440 669866 471822 669882
rect 476500 669868 476528 672590
rect 490564 672512 490616 672518
rect 490564 672454 490616 672460
rect 518714 672480 518770 672489
rect 481180 671084 481232 671090
rect 481180 671026 481232 671032
rect 481192 669868 481220 671026
rect 485792 669866 485898 669882
rect 490576 669868 490604 672454
rect 518714 672415 518770 672424
rect 499948 672172 500000 672178
rect 499948 672114 500000 672120
rect 500868 672172 500920 672178
rect 500868 672114 500920 672120
rect 495256 670948 495308 670954
rect 495256 670890 495308 670896
rect 495268 669868 495296 670890
rect 499960 669868 499988 672114
rect 500880 669866 500908 672114
rect 504640 672104 504692 672110
rect 504640 672046 504692 672052
rect 504652 669868 504680 672046
rect 509332 670880 509384 670886
rect 509332 670822 509384 670828
rect 509344 669868 509372 670822
rect 513760 669866 514050 669882
rect 518728 669868 518756 672415
rect 532790 672344 532846 672353
rect 532790 672279 532846 672288
rect 523406 670984 523462 670993
rect 523406 670919 523462 670928
rect 523420 669868 523448 670919
rect 527744 669866 528126 669882
rect 532804 669868 532832 672279
rect 546866 672208 546922 672217
rect 542176 672172 542228 672178
rect 546866 672143 546922 672152
rect 542176 672114 542228 672120
rect 537482 670848 537538 670857
rect 537482 670783 537538 670792
rect 537496 669868 537524 670783
rect 542188 669868 542216 672114
rect 546880 669868 546908 672143
rect 554044 671628 554096 671634
rect 554044 671570 554096 671576
rect 443276 669860 443578 669866
rect 429200 669802 429252 669808
rect 443328 669854 443578 669860
rect 457444 669860 457746 669866
rect 443276 669802 443328 669808
rect 457496 669854 457746 669860
rect 471428 669860 471822 669866
rect 457444 669802 457496 669808
rect 471480 669854 471822 669860
rect 485780 669860 485898 669866
rect 471428 669802 471480 669808
rect 485832 669854 485898 669860
rect 500868 669860 500920 669866
rect 485780 669802 485832 669808
rect 500868 669802 500920 669808
rect 513748 669860 514050 669866
rect 513800 669854 514050 669860
rect 527732 669860 528126 669866
rect 513748 669802 513800 669808
rect 527784 669854 528126 669860
rect 527732 669802 527784 669808
rect 133880 669792 133932 669798
rect 129030 669730 129320 669746
rect 133722 669740 133880 669746
rect 152832 669792 152884 669798
rect 133722 669734 133932 669740
rect 152490 669740 152832 669746
rect 152490 669734 152884 669740
rect 129030 669724 129332 669730
rect 129030 669718 129280 669724
rect 133722 669718 133920 669734
rect 152490 669718 152872 669734
rect 129280 669666 129332 669672
rect 110328 669656 110380 669662
rect 30654 669624 30710 669633
rect 30406 669582 30654 669610
rect 100786 669594 101168 669610
rect 110170 669604 110328 669610
rect 110170 669598 110380 669604
rect 100786 669588 101180 669594
rect 100786 669582 101128 669588
rect 30654 669559 30710 669568
rect 110170 669582 110368 669598
rect 101128 669530 101180 669536
rect 63408 669520 63460 669526
rect 16486 669488 16542 669497
rect 16330 669446 16486 669474
rect 21270 669488 21326 669497
rect 21022 669446 21270 669474
rect 16486 669423 16542 669432
rect 25714 669446 26004 669474
rect 39790 669458 39988 669474
rect 39790 669452 40000 669458
rect 39790 669446 39948 669452
rect 21270 669423 21326 669432
rect 25976 669390 26004 669446
rect 49174 669446 49464 669474
rect 53866 669446 54248 669474
rect 63250 669468 63408 669474
rect 72976 669520 73028 669526
rect 63250 669462 63460 669468
rect 72634 669468 72976 669474
rect 72634 669462 73028 669468
rect 63250 669446 63448 669462
rect 72634 669446 73016 669462
rect 39948 669394 40000 669400
rect 49436 669390 49464 669446
rect 54220 669390 54248 669446
rect 25964 669384 26016 669390
rect 25964 669326 26016 669332
rect 49424 669384 49476 669390
rect 49424 669326 49476 669332
rect 54208 669384 54260 669390
rect 54208 669326 54260 669332
rect 194704 669254 194732 669324
rect 194692 669248 194744 669254
rect 194692 669190 194744 669196
rect 13452 502308 13504 502314
rect 13452 502250 13504 502256
rect 554056 485790 554084 671570
rect 555424 671016 555476 671022
rect 555424 670958 555476 670964
rect 554136 668908 554188 668914
rect 554136 668850 554188 668856
rect 554148 578202 554176 668850
rect 554136 578196 554188 578202
rect 554136 578138 554188 578144
rect 554044 485784 554096 485790
rect 554044 485726 554096 485732
rect 13360 423632 13412 423638
rect 13360 423574 13412 423580
rect 555436 206990 555464 670958
rect 555528 525774 555556 673202
rect 566648 673056 566700 673062
rect 566648 672998 566700 673004
rect 558276 672444 558328 672450
rect 558276 672386 558328 672392
rect 556988 671764 557040 671770
rect 556988 671706 557040 671712
rect 555608 670132 555660 670138
rect 555608 670074 555660 670080
rect 555620 538218 555648 670074
rect 556802 669352 556858 669361
rect 556802 669287 556858 669296
rect 555608 538212 555660 538218
rect 555608 538154 555660 538160
rect 555516 525768 555568 525774
rect 555516 525710 555568 525716
rect 555424 206984 555476 206990
rect 555424 206926 555476 206932
rect 13268 202836 13320 202842
rect 13268 202778 13320 202784
rect 13176 164212 13228 164218
rect 13176 164154 13228 164160
rect 13084 59356 13136 59362
rect 13084 59298 13136 59304
rect 12256 48272 12308 48278
rect 12256 48214 12308 48220
rect 10968 47524 11020 47530
rect 10968 47466 11020 47472
rect 10324 20664 10376 20670
rect 10324 20606 10376 20612
rect 10980 3534 11008 47466
rect 12268 3534 12296 48214
rect 12348 48068 12400 48074
rect 12348 48010 12400 48016
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 7668 480 7696 3470
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 12360 480 12388 48010
rect 13728 48000 13780 48006
rect 13728 47942 13780 47948
rect 13740 6914 13768 47942
rect 14476 47598 14504 50116
rect 15488 47802 15516 50116
rect 16592 48210 16620 50116
rect 16580 48204 16632 48210
rect 16580 48146 16632 48152
rect 15476 47796 15528 47802
rect 15476 47738 15528 47744
rect 17696 47666 17724 50116
rect 17868 48204 17920 48210
rect 17868 48146 17920 48152
rect 17684 47660 17736 47666
rect 17684 47602 17736 47608
rect 14464 47592 14516 47598
rect 14464 47534 14516 47540
rect 15108 47456 15160 47462
rect 15108 47398 15160 47404
rect 15120 6914 15148 47398
rect 16488 47388 16540 47394
rect 16488 47330 16540 47336
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3534 16528 47330
rect 17880 3534 17908 48146
rect 18800 47870 18828 50116
rect 19904 47938 19932 50116
rect 21008 48142 21036 50116
rect 20996 48136 21048 48142
rect 20996 48078 21048 48084
rect 19892 47932 19944 47938
rect 19892 47874 19944 47880
rect 18788 47864 18840 47870
rect 18788 47806 18840 47812
rect 19248 47864 19300 47870
rect 19248 47806 19300 47812
rect 19260 3534 19288 47806
rect 20628 47796 20680 47802
rect 20628 47738 20680 47744
rect 20536 47592 20588 47598
rect 20536 47534 20588 47540
rect 20548 16574 20576 47534
rect 20456 16546 20576 16574
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 15948 480 15976 3470
rect 17052 480 17080 3470
rect 18248 480 18276 3470
rect 19444 480 19472 3538
rect 20456 3482 20484 16546
rect 20640 6914 20668 47738
rect 22112 47734 22140 50116
rect 22100 47728 22152 47734
rect 22100 47670 22152 47676
rect 23216 47530 23244 50116
rect 24320 48278 24348 50116
rect 24308 48272 24360 48278
rect 24308 48214 24360 48220
rect 24768 48136 24820 48142
rect 24768 48078 24820 48084
rect 23388 47728 23440 47734
rect 23388 47670 23440 47676
rect 23204 47524 23256 47530
rect 23204 47466 23256 47472
rect 22008 47320 22060 47326
rect 22008 47262 22060 47268
rect 22020 6914 22048 47262
rect 23400 6914 23428 47670
rect 20548 6886 20668 6914
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20548 3602 20576 6886
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 20456 3454 20668 3482
rect 20640 480 20668 3454
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3534 24808 48078
rect 25424 48074 25452 50116
rect 25412 48068 25464 48074
rect 25412 48010 25464 48016
rect 26436 48006 26464 50116
rect 27436 48272 27488 48278
rect 27436 48214 27488 48220
rect 26424 48000 26476 48006
rect 26424 47942 26476 47948
rect 26148 47932 26200 47938
rect 26148 47874 26200 47880
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24228 480 24256 3470
rect 26160 2990 26188 47874
rect 27448 45554 27476 48214
rect 27540 47462 27568 50116
rect 27528 47456 27580 47462
rect 27528 47398 27580 47404
rect 28644 47394 28672 50116
rect 29748 48210 29776 50116
rect 29736 48204 29788 48210
rect 29736 48146 29788 48152
rect 28908 48068 28960 48074
rect 28908 48010 28960 48016
rect 28816 47660 28868 47666
rect 28816 47602 28868 47608
rect 28632 47388 28684 47394
rect 28632 47330 28684 47336
rect 27448 45526 27568 45554
rect 27540 3534 27568 45526
rect 28828 16574 28856 47602
rect 28736 16546 28856 16574
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 26148 2984 26200 2990
rect 26148 2926 26200 2932
rect 25332 480 25360 2926
rect 26528 480 26556 3470
rect 27724 480 27752 3538
rect 28736 3482 28764 16546
rect 28920 6914 28948 48010
rect 30288 48000 30340 48006
rect 30288 47942 30340 47948
rect 30300 6914 30328 47942
rect 30852 47870 30880 50116
rect 30840 47864 30892 47870
rect 30840 47806 30892 47812
rect 31668 47864 31720 47870
rect 31668 47806 31720 47812
rect 31680 6914 31708 47806
rect 31956 47802 31984 50116
rect 32784 50102 33074 50130
rect 31944 47796 31996 47802
rect 31944 47738 31996 47744
rect 32784 47598 32812 50102
rect 33048 48204 33100 48210
rect 33048 48146 33100 48152
rect 32772 47592 32824 47598
rect 32772 47534 32824 47540
rect 28828 6886 28948 6914
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 28828 3602 28856 6886
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 28736 3454 28948 3482
rect 28920 480 28948 3454
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 33060 3534 33088 48146
rect 34164 47326 34192 50116
rect 35268 47734 35296 50116
rect 36372 48142 36400 50116
rect 36360 48136 36412 48142
rect 36360 48078 36412 48084
rect 37476 47938 37504 50116
rect 38488 48278 38516 50116
rect 38476 48272 38528 48278
rect 38476 48214 38528 48220
rect 39592 48074 39620 50116
rect 39580 48068 39632 48074
rect 39580 48010 39632 48016
rect 39948 48068 40000 48074
rect 39948 48010 40000 48016
rect 37464 47932 37516 47938
rect 37464 47874 37516 47880
rect 38568 47932 38620 47938
rect 38568 47874 38620 47880
rect 35808 47796 35860 47802
rect 35808 47738 35860 47744
rect 35256 47728 35308 47734
rect 35256 47670 35308 47676
rect 34428 47524 34480 47530
rect 34428 47466 34480 47472
rect 34152 47320 34204 47326
rect 34152 47262 34204 47268
rect 34440 3534 34468 47466
rect 35820 3534 35848 47738
rect 37096 47728 37148 47734
rect 37096 47670 37148 47676
rect 37108 3534 37136 47670
rect 37188 47592 37240 47598
rect 37188 47534 37240 47540
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 34808 480 34836 3470
rect 36004 480 36032 3470
rect 37200 480 37228 47534
rect 38580 6914 38608 47874
rect 39960 6914 39988 48010
rect 40696 47666 40724 50116
rect 41328 48136 41380 48142
rect 41328 48078 41380 48084
rect 40684 47660 40736 47666
rect 40684 47602 40736 47608
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3534 41368 48078
rect 41800 48006 41828 50116
rect 41788 48000 41840 48006
rect 41788 47942 41840 47948
rect 42708 48000 42760 48006
rect 42708 47942 42760 47948
rect 42720 3534 42748 47942
rect 42904 47870 42932 50116
rect 44008 48210 44036 50116
rect 43996 48204 44048 48210
rect 43996 48146 44048 48152
rect 42892 47864 42944 47870
rect 42892 47806 42944 47812
rect 44088 47864 44140 47870
rect 44088 47806 44140 47812
rect 44100 3534 44128 47806
rect 45112 47530 45140 50116
rect 45468 48272 45520 48278
rect 45468 48214 45520 48220
rect 45376 47660 45428 47666
rect 45376 47602 45428 47608
rect 45100 47524 45152 47530
rect 45100 47466 45152 47472
rect 45388 16574 45416 47602
rect 45296 16546 45416 16574
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 3538
rect 45296 3482 45324 16546
rect 45480 6914 45508 48214
rect 46216 47802 46244 50116
rect 46204 47796 46256 47802
rect 46204 47738 46256 47744
rect 46848 47796 46900 47802
rect 46848 47738 46900 47744
rect 46860 6914 46888 47738
rect 47320 47734 47348 50116
rect 48228 48204 48280 48210
rect 48228 48146 48280 48152
rect 47308 47728 47360 47734
rect 47308 47670 47360 47676
rect 48240 6914 48268 48146
rect 48424 47598 48452 50116
rect 49528 47938 49556 50116
rect 50540 48074 50568 50116
rect 51644 48142 51672 50116
rect 51632 48136 51684 48142
rect 51632 48078 51684 48084
rect 52368 48136 52420 48142
rect 52368 48078 52420 48084
rect 50528 48068 50580 48074
rect 50528 48010 50580 48016
rect 50988 48068 51040 48074
rect 50988 48010 51040 48016
rect 49516 47932 49568 47938
rect 49516 47874 49568 47880
rect 48412 47592 48464 47598
rect 48412 47534 48464 47540
rect 49608 47592 49660 47598
rect 49608 47534 49660 47540
rect 45388 6886 45508 6914
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 45388 3602 45416 6886
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45296 3454 45508 3482
rect 45480 480 45508 3454
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3534 49648 47534
rect 51000 3534 51028 48010
rect 52380 3534 52408 48078
rect 52748 48006 52776 50116
rect 52736 48000 52788 48006
rect 52736 47942 52788 47948
rect 53656 47932 53708 47938
rect 53656 47874 53708 47880
rect 53668 3534 53696 47874
rect 53852 47870 53880 50116
rect 54956 48278 54984 50116
rect 54944 48272 54996 48278
rect 54944 48214 54996 48220
rect 53840 47864 53892 47870
rect 53840 47806 53892 47812
rect 55128 47864 55180 47870
rect 55128 47806 55180 47812
rect 53748 47728 53800 47734
rect 53748 47670 53800 47676
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 53656 3528 53708 3534
rect 53656 3470 53708 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51368 480 51396 3470
rect 52564 480 52592 3470
rect 53760 480 53788 47670
rect 55140 6914 55168 47806
rect 56060 47666 56088 50116
rect 57164 47802 57192 50116
rect 58268 48210 58296 50116
rect 58256 48204 58308 48210
rect 58256 48146 58308 48152
rect 59268 48204 59320 48210
rect 59268 48146 59320 48152
rect 57152 47796 57204 47802
rect 57152 47738 57204 47744
rect 57888 47796 57940 47802
rect 57888 47738 57940 47744
rect 56048 47660 56100 47666
rect 56048 47602 56100 47608
rect 56508 47660 56560 47666
rect 56508 47602 56560 47608
rect 54956 6886 55168 6914
rect 54956 480 54984 6886
rect 56520 3534 56548 47602
rect 57900 3534 57928 47738
rect 59280 3534 59308 48146
rect 59372 47598 59400 50116
rect 60476 48074 60504 50116
rect 61488 48142 61516 50116
rect 61476 48136 61528 48142
rect 61476 48078 61528 48084
rect 60464 48068 60516 48074
rect 60464 48010 60516 48016
rect 61936 48068 61988 48074
rect 61936 48010 61988 48016
rect 59360 47592 59412 47598
rect 59360 47534 59412 47540
rect 60648 47592 60700 47598
rect 60648 47534 60700 47540
rect 60660 3534 60688 47534
rect 61948 3534 61976 48010
rect 62028 48000 62080 48006
rect 62028 47942 62080 47948
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56508 3528 56560 3534
rect 56508 3470 56560 3476
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 60832 3528 60884 3534
rect 60832 3470 60884 3476
rect 61936 3528 61988 3534
rect 61936 3470 61988 3476
rect 56060 480 56088 3470
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 59648 480 59676 3470
rect 60844 480 60872 3470
rect 62040 480 62068 47942
rect 62592 47938 62620 50116
rect 62580 47932 62632 47938
rect 62580 47874 62632 47880
rect 63408 47932 63460 47938
rect 63408 47874 63460 47880
rect 63420 6914 63448 47874
rect 63696 47734 63724 50116
rect 64800 47870 64828 50116
rect 64788 47864 64840 47870
rect 64788 47806 64840 47812
rect 63684 47728 63736 47734
rect 63684 47670 63736 47676
rect 64788 47728 64840 47734
rect 64788 47670 64840 47676
rect 63236 6886 63448 6914
rect 63236 480 63264 6886
rect 64800 3534 64828 47670
rect 65904 47666 65932 50116
rect 67008 47802 67036 50116
rect 68112 48210 68140 50116
rect 68100 48204 68152 48210
rect 68100 48146 68152 48152
rect 67548 48136 67600 48142
rect 67548 48078 67600 48084
rect 66996 47796 67048 47802
rect 66996 47738 67048 47744
rect 66168 47728 66220 47734
rect 66168 47670 66220 47676
rect 65892 47660 65944 47666
rect 65892 47602 65944 47608
rect 66180 3534 66208 47670
rect 67560 3534 67588 48078
rect 69216 47598 69244 50116
rect 70320 48074 70348 50116
rect 70308 48068 70360 48074
rect 70308 48010 70360 48016
rect 71424 48006 71452 50116
rect 71412 48000 71464 48006
rect 71412 47942 71464 47948
rect 70308 47932 70360 47938
rect 70308 47874 70360 47880
rect 69204 47592 69256 47598
rect 69204 47534 69256 47540
rect 70216 47592 70268 47598
rect 70216 47534 70268 47540
rect 68928 46980 68980 46986
rect 68928 46922 68980 46928
rect 68940 3534 68968 46922
rect 70228 16574 70256 47534
rect 70136 16546 70256 16574
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 64328 3528 64380 3534
rect 64328 3470 64380 3476
rect 64788 3528 64840 3534
rect 64788 3470 64840 3476
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 66720 3528 66772 3534
rect 66720 3470 66772 3476
rect 67548 3528 67600 3534
rect 67548 3470 67600 3476
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 64340 480 64368 3470
rect 65536 480 65564 3470
rect 66732 480 66760 3470
rect 67928 480 67956 3470
rect 69124 480 69152 3538
rect 70136 3482 70164 16546
rect 70320 6914 70348 47874
rect 72528 47870 72556 50116
rect 73068 48204 73120 48210
rect 73068 48146 73120 48152
rect 72516 47864 72568 47870
rect 72516 47806 72568 47812
rect 71688 47660 71740 47666
rect 71688 47602 71740 47608
rect 71700 6914 71728 47602
rect 70228 6886 70348 6914
rect 71516 6886 71728 6914
rect 70228 3602 70256 6886
rect 70216 3596 70268 3602
rect 70216 3538 70268 3544
rect 70136 3454 70348 3482
rect 70320 480 70348 3454
rect 71516 480 71544 6886
rect 73080 3534 73108 48146
rect 73540 47530 73568 50116
rect 74448 47932 74500 47938
rect 74448 47874 74500 47880
rect 73528 47524 73580 47530
rect 73528 47466 73580 47472
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 72620 480 72648 3470
rect 74460 3466 74488 47874
rect 74644 47870 74672 50116
rect 75748 48142 75776 50116
rect 75736 48136 75788 48142
rect 75736 48078 75788 48084
rect 74632 47864 74684 47870
rect 74632 47806 74684 47812
rect 75828 47456 75880 47462
rect 75828 47398 75880 47404
rect 75840 3534 75868 47398
rect 76852 46986 76880 50116
rect 77956 48074 77984 50116
rect 77944 48068 77996 48074
rect 77944 48010 77996 48016
rect 77208 47796 77260 47802
rect 77208 47738 77260 47744
rect 76840 46980 76892 46986
rect 76840 46922 76892 46928
rect 77220 3534 77248 47738
rect 79060 47598 79088 50116
rect 79968 48068 80020 48074
rect 79968 48010 80020 48016
rect 79048 47592 79100 47598
rect 79048 47534 79100 47540
rect 78496 47048 78548 47054
rect 78496 46990 78548 46996
rect 78508 16574 78536 46990
rect 78588 46980 78640 46986
rect 78588 46922 78640 46928
rect 78416 16546 78536 16574
rect 77392 3596 77444 3602
rect 77392 3538 77444 3544
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 73804 3460 73856 3466
rect 73804 3402 73856 3408
rect 74448 3460 74500 3466
rect 74448 3402 74500 3408
rect 73816 480 73844 3402
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77404 480 77432 3538
rect 78416 3482 78444 16546
rect 78600 6914 78628 46922
rect 79980 6914 80008 48010
rect 80164 47666 80192 50116
rect 81268 48210 81296 50116
rect 81256 48204 81308 48210
rect 81256 48146 81308 48152
rect 82372 47938 82400 50116
rect 82360 47932 82412 47938
rect 82360 47874 82412 47880
rect 80152 47660 80204 47666
rect 80152 47602 80204 47608
rect 81348 47660 81400 47666
rect 81348 47602 81400 47608
rect 78508 6886 78628 6914
rect 79704 6886 80008 6914
rect 78508 3602 78536 6886
rect 78496 3596 78548 3602
rect 78496 3538 78548 3544
rect 78416 3454 78628 3482
rect 78600 480 78628 3454
rect 79704 480 79732 6886
rect 81360 3330 81388 47602
rect 82728 47592 82780 47598
rect 82728 47534 82780 47540
rect 82740 3534 82768 47534
rect 83476 47462 83504 50116
rect 84108 47864 84160 47870
rect 84108 47806 84160 47812
rect 83464 47456 83516 47462
rect 83464 47398 83516 47404
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 82728 3528 82780 3534
rect 82728 3470 82780 3476
rect 80888 3324 80940 3330
rect 80888 3266 80940 3272
rect 81348 3324 81400 3330
rect 81348 3266 81400 3272
rect 80900 480 80928 3266
rect 82096 480 82124 3470
rect 84120 2990 84148 47806
rect 84580 47802 84608 50116
rect 84568 47796 84620 47802
rect 84568 47738 84620 47744
rect 85488 47728 85540 47734
rect 85488 47670 85540 47676
rect 85500 3262 85528 47670
rect 85592 46986 85620 50116
rect 86696 47054 86724 50116
rect 87800 48074 87828 50116
rect 87788 48068 87840 48074
rect 87788 48010 87840 48016
rect 86776 47932 86828 47938
rect 86776 47874 86828 47880
rect 86684 47048 86736 47054
rect 86684 46990 86736 46996
rect 85580 46980 85632 46986
rect 85580 46922 85632 46928
rect 86788 3330 86816 47874
rect 86868 47796 86920 47802
rect 86868 47738 86920 47744
rect 85672 3324 85724 3330
rect 85672 3266 85724 3272
rect 86776 3324 86828 3330
rect 86776 3266 86828 3272
rect 84476 3256 84528 3262
rect 84476 3198 84528 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 83280 2984 83332 2990
rect 83280 2926 83332 2932
rect 84108 2984 84160 2990
rect 84108 2926 84160 2932
rect 83292 480 83320 2926
rect 84488 480 84516 3198
rect 85684 480 85712 3266
rect 86880 480 86908 47738
rect 88904 47666 88932 50116
rect 88892 47660 88944 47666
rect 88892 47602 88944 47608
rect 89628 47660 89680 47666
rect 89628 47602 89680 47608
rect 88248 46980 88300 46986
rect 88248 46922 88300 46928
rect 88260 6914 88288 46922
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 89640 3330 89668 47602
rect 90008 47598 90036 50116
rect 91008 48068 91060 48074
rect 91008 48010 91060 48016
rect 89996 47592 90048 47598
rect 89996 47534 90048 47540
rect 91020 3534 91048 48010
rect 91112 47870 91140 50116
rect 91100 47864 91152 47870
rect 91100 47806 91152 47812
rect 92216 47734 92244 50116
rect 92388 48000 92440 48006
rect 92388 47942 92440 47948
rect 92204 47728 92256 47734
rect 92204 47670 92256 47676
rect 92400 3534 92428 47942
rect 93320 47938 93348 50116
rect 93308 47932 93360 47938
rect 93308 47874 93360 47880
rect 93768 47864 93820 47870
rect 93768 47806 93820 47812
rect 93780 3534 93808 47806
rect 94424 47802 94452 50116
rect 95056 48136 95108 48142
rect 95056 48078 95108 48084
rect 94412 47796 94464 47802
rect 94412 47738 94464 47744
rect 95068 16574 95096 48078
rect 95148 47320 95200 47326
rect 95148 47262 95200 47268
rect 94976 16546 95096 16574
rect 93952 3596 94004 3602
rect 93952 3538 94004 3544
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 92388 3528 92440 3534
rect 92388 3470 92440 3476
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 89168 3324 89220 3330
rect 89168 3266 89220 3272
rect 89628 3324 89680 3330
rect 89628 3266 89680 3272
rect 89180 480 89208 3266
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 92768 480 92796 3470
rect 93964 480 93992 3538
rect 94976 3482 95004 16546
rect 95160 6914 95188 47262
rect 95528 46986 95556 50116
rect 96632 47666 96660 50116
rect 97644 48074 97672 50116
rect 97632 48068 97684 48074
rect 97632 48010 97684 48016
rect 98748 48006 98776 50116
rect 98736 48000 98788 48006
rect 98736 47942 98788 47948
rect 99852 47870 99880 50116
rect 99840 47864 99892 47870
rect 99840 47806 99892 47812
rect 100668 47796 100720 47802
rect 100668 47738 100720 47744
rect 96620 47660 96672 47666
rect 96620 47602 96672 47608
rect 96528 47456 96580 47462
rect 96528 47398 96580 47404
rect 95516 46980 95568 46986
rect 95516 46922 95568 46928
rect 96540 6914 96568 47398
rect 99288 47048 99340 47054
rect 99288 46990 99340 46996
rect 97908 46980 97960 46986
rect 97908 46922 97960 46928
rect 95068 6886 95188 6914
rect 96264 6886 96568 6914
rect 95068 3602 95096 6886
rect 95056 3596 95108 3602
rect 95056 3538 95108 3544
rect 94976 3454 95188 3482
rect 95160 480 95188 3454
rect 96264 480 96292 6886
rect 97920 3534 97948 46922
rect 99300 3534 99328 46990
rect 100680 3534 100708 47738
rect 100956 47326 100984 50116
rect 102060 48142 102088 50116
rect 102048 48136 102100 48142
rect 102048 48078 102100 48084
rect 102048 48000 102100 48006
rect 102048 47942 102100 47948
rect 100944 47320 100996 47326
rect 100944 47262 100996 47268
rect 102060 3534 102088 47942
rect 103164 47462 103192 50116
rect 103336 47932 103388 47938
rect 103336 47874 103388 47880
rect 103152 47456 103204 47462
rect 103152 47398 103204 47404
rect 103348 16574 103376 47874
rect 103428 47728 103480 47734
rect 103428 47670 103480 47676
rect 103256 16546 103376 16574
rect 103256 3534 103284 16546
rect 103440 6914 103468 47670
rect 104268 46986 104296 50116
rect 104808 47660 104860 47666
rect 104808 47602 104860 47608
rect 104256 46980 104308 46986
rect 104256 46922 104308 46928
rect 104820 6914 104848 47602
rect 105372 47054 105400 50116
rect 106476 47802 106504 50116
rect 107580 48006 107608 50116
rect 107568 48000 107620 48006
rect 107568 47942 107620 47948
rect 108592 47938 108620 50116
rect 108580 47932 108632 47938
rect 108580 47874 108632 47880
rect 107568 47864 107620 47870
rect 107568 47806 107620 47812
rect 106464 47796 106516 47802
rect 106464 47738 106516 47744
rect 106188 47592 106240 47598
rect 106188 47534 106240 47540
rect 105360 47048 105412 47054
rect 105360 46990 105412 46996
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 102232 3528 102284 3534
rect 102232 3470 102284 3476
rect 103244 3528 103296 3534
rect 103244 3470 103296 3476
rect 97460 480 97488 3470
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 101048 480 101076 3470
rect 102244 480 102272 3470
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 106200 3534 106228 47534
rect 107580 3534 107608 47806
rect 109696 47734 109724 50116
rect 109684 47728 109736 47734
rect 109684 47670 109736 47676
rect 110800 47666 110828 50116
rect 111616 47728 111668 47734
rect 111616 47670 111668 47676
rect 110788 47660 110840 47666
rect 110788 47602 110840 47608
rect 110328 47116 110380 47122
rect 110328 47058 110380 47064
rect 108948 47048 109000 47054
rect 108948 46990 109000 46996
rect 108960 3534 108988 46990
rect 110340 3534 110368 47058
rect 111628 16574 111656 47670
rect 111708 47660 111760 47666
rect 111708 47602 111760 47608
rect 111536 16546 111656 16574
rect 111536 3534 111564 16546
rect 111720 6914 111748 47602
rect 111904 47598 111932 50116
rect 113008 47870 113036 50116
rect 112996 47864 113048 47870
rect 112996 47806 113048 47812
rect 113088 47796 113140 47802
rect 113088 47738 113140 47744
rect 111892 47592 111944 47598
rect 111892 47534 111944 47540
rect 113100 6914 113128 47738
rect 114112 47054 114140 50116
rect 114468 47864 114520 47870
rect 114468 47806 114520 47812
rect 114100 47048 114152 47054
rect 114100 46990 114152 46996
rect 111628 6886 111748 6914
rect 112824 6886 113128 6914
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 110328 3528 110380 3534
rect 110328 3470 110380 3476
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 111524 3528 111576 3534
rect 111524 3470 111576 3476
rect 105740 480 105768 3470
rect 106936 480 106964 3470
rect 108132 480 108160 3470
rect 109328 480 109356 3470
rect 110524 480 110552 3470
rect 111628 480 111656 6886
rect 112824 480 112852 6886
rect 114480 3534 114508 47806
rect 115216 47122 115244 50116
rect 115848 47932 115900 47938
rect 115848 47874 115900 47880
rect 115204 47116 115256 47122
rect 115204 47058 115256 47064
rect 115860 3534 115888 47874
rect 116320 47734 116348 50116
rect 116308 47728 116360 47734
rect 116308 47670 116360 47676
rect 117228 47728 117280 47734
rect 117228 47670 117280 47676
rect 117240 3534 117268 47670
rect 117424 47666 117452 50116
rect 118528 47802 118556 50116
rect 119632 47870 119660 50116
rect 120644 47938 120672 50116
rect 120632 47932 120684 47938
rect 120632 47874 120684 47880
rect 119620 47864 119672 47870
rect 119620 47806 119672 47812
rect 118516 47796 118568 47802
rect 118516 47738 118568 47744
rect 121368 47796 121420 47802
rect 121368 47738 121420 47744
rect 117412 47660 117464 47666
rect 117412 47602 117464 47608
rect 119896 47184 119948 47190
rect 119896 47126 119948 47132
rect 118608 47048 118660 47054
rect 118608 46990 118660 46996
rect 118620 3534 118648 46990
rect 114008 3528 114060 3534
rect 114008 3470 114060 3476
rect 114468 3528 114520 3534
rect 114468 3470 114520 3476
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 117228 3528 117280 3534
rect 117228 3470 117280 3476
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 118608 3528 118660 3534
rect 118608 3470 118660 3476
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 114020 480 114048 3470
rect 115216 480 115244 3470
rect 116412 480 116440 3470
rect 117608 480 117636 3470
rect 118804 480 118832 3470
rect 119908 480 119936 47126
rect 119988 46980 120040 46986
rect 119988 46922 120040 46928
rect 120000 3534 120028 46922
rect 121380 6914 121408 47738
rect 121748 47734 121776 50116
rect 121736 47728 121788 47734
rect 121736 47670 121788 47676
rect 122748 47728 122800 47734
rect 122748 47670 122800 47676
rect 121104 6886 121408 6914
rect 119988 3528 120040 3534
rect 119988 3470 120040 3476
rect 121104 480 121132 6886
rect 122760 3534 122788 47670
rect 122852 47054 122880 50116
rect 122840 47048 122892 47054
rect 122840 46990 122892 46996
rect 123956 46986 123984 50116
rect 124128 47320 124180 47326
rect 124128 47262 124180 47268
rect 123944 46980 123996 46986
rect 123944 46922 123996 46928
rect 124140 3534 124168 47262
rect 125060 47190 125088 50116
rect 126164 47802 126192 50116
rect 126152 47796 126204 47802
rect 126152 47738 126204 47744
rect 126888 47796 126940 47802
rect 126888 47738 126940 47744
rect 125048 47184 125100 47190
rect 125048 47126 125100 47132
rect 125508 47048 125560 47054
rect 125508 46990 125560 46996
rect 125520 3534 125548 46990
rect 126900 3534 126928 47738
rect 127268 47734 127296 50116
rect 127256 47728 127308 47734
rect 127256 47670 127308 47676
rect 128372 47326 128400 50116
rect 128360 47320 128412 47326
rect 128360 47262 128412 47268
rect 128268 47184 128320 47190
rect 128268 47126 128320 47132
rect 128280 6914 128308 47126
rect 129476 47054 129504 50116
rect 130384 47864 130436 47870
rect 130384 47806 130436 47812
rect 129464 47048 129516 47054
rect 129464 46990 129516 46996
rect 129648 47048 129700 47054
rect 129648 46990 129700 46996
rect 129660 6914 129688 46990
rect 128188 6886 128308 6914
rect 129384 6886 129688 6914
rect 122288 3528 122340 3534
rect 122288 3470 122340 3476
rect 122748 3528 122800 3534
rect 122748 3470 122800 3476
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 126888 3528 126940 3534
rect 126888 3470 126940 3476
rect 122300 480 122328 3470
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125888 480 125916 3470
rect 126980 3324 127032 3330
rect 126980 3266 127032 3272
rect 126992 480 127020 3266
rect 128188 480 128216 6886
rect 129384 480 129412 6886
rect 130396 3330 130424 47806
rect 130580 47802 130608 50116
rect 131684 47870 131712 50116
rect 131672 47864 131724 47870
rect 131672 47806 131724 47812
rect 130568 47796 130620 47802
rect 130568 47738 130620 47744
rect 132408 47796 132460 47802
rect 132408 47738 132460 47744
rect 131028 47116 131080 47122
rect 131028 47058 131080 47064
rect 131040 3534 131068 47058
rect 130568 3528 130620 3534
rect 130568 3470 130620 3476
rect 131028 3528 131080 3534
rect 131028 3470 131080 3476
rect 130384 3324 130436 3330
rect 130384 3266 130436 3272
rect 130580 480 130608 3470
rect 132420 3466 132448 47738
rect 132696 47190 132724 50116
rect 132684 47184 132736 47190
rect 132684 47126 132736 47132
rect 133800 47054 133828 50116
rect 134904 47122 134932 50116
rect 135168 47932 135220 47938
rect 135168 47874 135220 47880
rect 134892 47116 134944 47122
rect 134892 47058 134944 47064
rect 133788 47048 133840 47054
rect 133788 46990 133840 46996
rect 133788 46912 133840 46918
rect 133788 46854 133840 46860
rect 133800 3534 133828 46854
rect 135180 3534 135208 47874
rect 136008 47802 136036 50116
rect 135996 47796 136048 47802
rect 135996 47738 136048 47744
rect 136548 47796 136600 47802
rect 136548 47738 136600 47744
rect 132960 3528 133012 3534
rect 132960 3470 133012 3476
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 134156 3528 134208 3534
rect 134156 3470 134208 3476
rect 135168 3528 135220 3534
rect 135168 3470 135220 3476
rect 136456 3528 136508 3534
rect 136456 3470 136508 3476
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 132408 3460 132460 3466
rect 132408 3402 132460 3408
rect 131776 480 131804 3402
rect 132972 480 133000 3470
rect 134168 480 134196 3470
rect 135260 3460 135312 3466
rect 135260 3402 135312 3408
rect 135272 480 135300 3402
rect 136468 480 136496 3470
rect 136560 3466 136588 47738
rect 137112 46986 137140 50116
rect 138216 47938 138244 50116
rect 138204 47932 138256 47938
rect 138204 47874 138256 47880
rect 137284 47864 137336 47870
rect 137284 47806 137336 47812
rect 137100 46980 137152 46986
rect 137100 46922 137152 46928
rect 137296 3534 137324 47806
rect 139320 47802 139348 50116
rect 140424 47870 140452 50116
rect 140412 47864 140464 47870
rect 140412 47806 140464 47812
rect 139308 47796 139360 47802
rect 139308 47738 139360 47744
rect 141528 47734 141556 50116
rect 137928 47728 137980 47734
rect 137928 47670 137980 47676
rect 141516 47728 141568 47734
rect 141516 47670 141568 47676
rect 137940 6914 137968 47670
rect 142632 47122 142660 50116
rect 143448 47456 143500 47462
rect 143448 47398 143500 47404
rect 139308 47116 139360 47122
rect 139308 47058 139360 47064
rect 142620 47116 142672 47122
rect 142620 47058 142672 47064
rect 137664 6886 137968 6914
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 136548 3460 136600 3466
rect 136548 3402 136600 3408
rect 137664 480 137692 6886
rect 139320 3534 139348 47058
rect 140688 47048 140740 47054
rect 140688 46990 140740 46996
rect 140700 3534 140728 46990
rect 142068 46980 142120 46986
rect 142068 46922 142120 46928
rect 142080 3534 142108 46922
rect 143460 3534 143488 47398
rect 143644 47054 143672 50116
rect 143632 47048 143684 47054
rect 143632 46990 143684 46996
rect 144748 46986 144776 50116
rect 144828 47864 144880 47870
rect 144828 47806 144880 47812
rect 144736 46980 144788 46986
rect 144736 46922 144788 46928
rect 144840 46866 144868 47806
rect 145852 47462 145880 50116
rect 146208 47932 146260 47938
rect 146208 47874 146260 47880
rect 145840 47456 145892 47462
rect 145840 47398 145892 47404
rect 144748 46838 144868 46866
rect 144748 16574 144776 46838
rect 144828 46776 144880 46782
rect 144828 46718 144880 46724
rect 144656 16546 144776 16574
rect 138848 3528 138900 3534
rect 138848 3470 138900 3476
rect 139308 3528 139360 3534
rect 139308 3470 139360 3476
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 140688 3528 140740 3534
rect 140688 3470 140740 3476
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 142068 3528 142120 3534
rect 142068 3470 142120 3476
rect 142436 3528 142488 3534
rect 142436 3470 142488 3476
rect 143448 3528 143500 3534
rect 143448 3470 143500 3476
rect 138860 480 138888 3470
rect 140056 480 140084 3470
rect 141252 480 141280 3470
rect 142448 480 142476 3470
rect 144656 3058 144684 16546
rect 144840 6914 144868 46718
rect 146220 6914 146248 47874
rect 146956 47870 146984 50116
rect 146944 47864 146996 47870
rect 146944 47806 146996 47812
rect 147588 47796 147640 47802
rect 147588 47738 147640 47744
rect 144748 6886 144868 6914
rect 145944 6886 146248 6914
rect 143540 3052 143592 3058
rect 143540 2994 143592 3000
rect 144644 3052 144696 3058
rect 144644 2994 144696 3000
rect 143552 480 143580 2994
rect 144748 480 144776 6886
rect 145944 480 145972 6886
rect 147600 3534 147628 47738
rect 148060 46986 148088 50116
rect 149164 47938 149192 50116
rect 149152 47932 149204 47938
rect 149152 47874 149204 47880
rect 148968 47864 149020 47870
rect 148968 47806 149020 47812
rect 148048 46980 148100 46986
rect 148048 46922 148100 46928
rect 148980 3534 149008 47806
rect 150268 47802 150296 50116
rect 151372 47870 151400 50116
rect 151360 47864 151412 47870
rect 151360 47806 151412 47812
rect 150256 47796 150308 47802
rect 150256 47738 150308 47744
rect 151728 47048 151780 47054
rect 151728 46990 151780 46996
rect 151084 46980 151136 46986
rect 151084 46922 151136 46928
rect 151096 3534 151124 46922
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 148324 3528 148376 3534
rect 148324 3470 148376 3476
rect 148968 3528 149020 3534
rect 148968 3470 149020 3476
rect 149520 3528 149572 3534
rect 149520 3470 149572 3476
rect 151084 3528 151136 3534
rect 151084 3470 151136 3476
rect 147140 480 147168 3470
rect 148336 480 148364 3470
rect 149532 480 149560 3470
rect 151740 3058 151768 46990
rect 152476 46986 152504 50116
rect 153108 47864 153160 47870
rect 153108 47806 153160 47812
rect 153016 47796 153068 47802
rect 153016 47738 153068 47744
rect 152464 46980 152516 46986
rect 152464 46922 152516 46928
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 150624 3052 150676 3058
rect 150624 2994 150676 3000
rect 151728 3052 151780 3058
rect 151728 2994 151780 3000
rect 150636 480 150664 2994
rect 151832 480 151860 3470
rect 153028 480 153056 47738
rect 153120 3534 153148 47806
rect 153580 47054 153608 50116
rect 154684 47870 154712 50116
rect 154672 47864 154724 47870
rect 154672 47806 154724 47812
rect 155696 47802 155724 50116
rect 156064 50102 156814 50130
rect 155868 47864 155920 47870
rect 155868 47806 155920 47812
rect 155684 47796 155736 47802
rect 155684 47738 155736 47744
rect 153568 47048 153620 47054
rect 153568 46990 153620 46996
rect 153108 3528 153160 3534
rect 153108 3470 153160 3476
rect 154212 3528 154264 3534
rect 154212 3470 154264 3476
rect 154224 480 154252 3470
rect 155880 3466 155908 47806
rect 156064 3534 156092 50102
rect 157904 47870 157932 50116
rect 158628 47932 158680 47938
rect 158628 47874 158680 47880
rect 157892 47864 157944 47870
rect 157892 47806 157944 47812
rect 157248 47660 157300 47666
rect 157248 47602 157300 47608
rect 157260 3534 157288 47602
rect 158640 3534 158668 47874
rect 159008 47666 159036 50116
rect 160112 47938 160140 50116
rect 160100 47932 160152 47938
rect 160100 47874 160152 47880
rect 161216 47870 161244 50116
rect 161584 50102 162334 50130
rect 161584 48328 161612 50102
rect 161446 48314 161612 48328
rect 161400 48300 161612 48314
rect 161400 48286 161474 48300
rect 160008 47864 160060 47870
rect 160008 47806 160060 47812
rect 161204 47864 161256 47870
rect 161204 47806 161256 47812
rect 158996 47660 159048 47666
rect 158996 47602 159048 47608
rect 160020 3534 160048 47806
rect 161296 46980 161348 46986
rect 161296 46922 161348 46928
rect 156052 3528 156104 3534
rect 156052 3470 156104 3476
rect 156604 3528 156656 3534
rect 156604 3470 156656 3476
rect 157248 3528 157300 3534
rect 157248 3470 157300 3476
rect 157800 3528 157852 3534
rect 157800 3470 157852 3476
rect 158628 3528 158680 3534
rect 158628 3470 158680 3476
rect 158904 3528 158956 3534
rect 158904 3470 158956 3476
rect 160008 3528 160060 3534
rect 160008 3470 160060 3476
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 155408 3460 155460 3466
rect 155408 3402 155460 3408
rect 155868 3460 155920 3466
rect 155868 3402 155920 3408
rect 155420 480 155448 3402
rect 156616 480 156644 3470
rect 157812 480 157840 3470
rect 158916 480 158944 3470
rect 160112 480 160140 3470
rect 161308 480 161336 46922
rect 161400 3534 161428 48286
rect 162768 47864 162820 47870
rect 162768 47806 162820 47812
rect 162780 6914 162808 47806
rect 163424 46986 163452 50116
rect 164528 47870 164556 50116
rect 164516 47864 164568 47870
rect 164516 47806 164568 47812
rect 165632 47666 165660 50116
rect 165724 50102 166750 50130
rect 164148 47660 164200 47666
rect 164148 47602 164200 47608
rect 165620 47660 165672 47666
rect 165620 47602 165672 47608
rect 163412 46980 163464 46986
rect 163412 46922 163464 46928
rect 162504 6886 162808 6914
rect 161388 3528 161440 3534
rect 161388 3470 161440 3476
rect 162504 480 162532 6886
rect 164160 3534 164188 47602
rect 165724 3534 165752 50102
rect 167748 47870 167776 50116
rect 168576 50102 168866 50130
rect 169772 50102 169970 50130
rect 170140 50102 171074 50130
rect 166908 47864 166960 47870
rect 166908 47806 166960 47812
rect 167736 47864 167788 47870
rect 167736 47806 167788 47812
rect 166920 3534 166948 47806
rect 168380 3596 168432 3602
rect 168380 3538 168432 3544
rect 163688 3528 163740 3534
rect 163688 3470 163740 3476
rect 164148 3528 164200 3534
rect 164148 3470 164200 3476
rect 164884 3528 164936 3534
rect 164884 3470 164936 3476
rect 165712 3528 165764 3534
rect 165712 3470 165764 3476
rect 166080 3528 166132 3534
rect 166080 3470 166132 3476
rect 166908 3528 166960 3534
rect 166908 3470 166960 3476
rect 167184 3528 167236 3534
rect 167184 3470 167236 3476
rect 163700 480 163728 3470
rect 164896 480 164924 3470
rect 166092 480 166120 3470
rect 167196 480 167224 3470
rect 168392 480 168420 3538
rect 168576 3534 168604 50102
rect 169772 47852 169800 50102
rect 169680 47824 169800 47852
rect 169680 3602 169708 47824
rect 170140 45554 170168 50102
rect 171140 48340 171192 48346
rect 169864 45526 170168 45554
rect 171060 48288 171140 48314
rect 171060 48286 171192 48288
rect 169864 6914 169892 45526
rect 171060 6914 171088 48286
rect 171140 48282 171192 48286
rect 172164 48278 172192 50116
rect 172624 50102 173282 50130
rect 173912 50102 174386 50130
rect 175292 50102 175490 50130
rect 175568 50102 176594 50130
rect 172152 48272 172204 48278
rect 172152 48214 172204 48220
rect 169772 6886 169892 6914
rect 170784 6886 171088 6914
rect 169668 3596 169720 3602
rect 169668 3538 169720 3544
rect 168564 3528 168616 3534
rect 169772 3482 169800 6886
rect 168564 3470 168616 3476
rect 169588 3454 169800 3482
rect 169588 480 169616 3454
rect 170784 480 170812 6886
rect 172624 3534 172652 50102
rect 173912 47818 173940 50102
rect 175292 47818 175320 50102
rect 173820 47790 173940 47818
rect 175200 47790 175320 47818
rect 173820 3534 173848 47790
rect 175200 3534 175228 47790
rect 175568 45554 175596 50102
rect 177684 47870 177712 50116
rect 178052 50102 178802 50130
rect 179524 50102 179814 50130
rect 180812 50102 180918 50130
rect 180996 50102 182022 50130
rect 182192 50102 183126 50130
rect 183572 50102 184230 50130
rect 184952 50102 185334 50130
rect 176660 47864 176712 47870
rect 176660 47806 176712 47812
rect 177672 47864 177724 47870
rect 177672 47806 177724 47812
rect 175384 45526 175596 45554
rect 175384 16574 175412 45526
rect 175384 16546 175504 16574
rect 171968 3528 172020 3534
rect 171968 3470 172020 3476
rect 172612 3528 172664 3534
rect 172612 3470 172664 3476
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 175188 3528 175240 3534
rect 175188 3470 175240 3476
rect 171980 480 172008 3470
rect 173176 480 173204 3470
rect 174280 480 174308 3470
rect 175476 480 175504 16546
rect 176672 480 176700 47806
rect 178052 3482 178080 50102
rect 179524 3534 179552 50102
rect 180812 48314 180840 50102
rect 180720 48286 180840 48314
rect 180720 3534 180748 48286
rect 180996 3534 181024 50102
rect 177868 3454 178080 3482
rect 179052 3528 179104 3534
rect 179052 3470 179104 3476
rect 179512 3528 179564 3534
rect 179512 3470 179564 3476
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 180984 3528 181036 3534
rect 180984 3470 181036 3476
rect 181444 3528 181496 3534
rect 181444 3470 181496 3476
rect 177868 480 177896 3454
rect 179064 480 179092 3470
rect 180260 480 180288 3470
rect 181456 480 181484 3470
rect 182192 490 182220 50102
rect 183572 16574 183600 50102
rect 183572 16546 183784 16574
rect 182376 598 182588 626
rect 182376 490 182404 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 462 182404 490
rect 182560 480 182588 598
rect 183756 480 183784 16546
rect 184952 480 184980 50102
rect 186320 47864 186372 47870
rect 186320 47806 186372 47812
rect 186332 3602 186360 47806
rect 186320 3596 186372 3602
rect 186320 3538 186372 3544
rect 186424 3482 186452 50116
rect 187528 47870 187556 50116
rect 187712 50102 188646 50130
rect 189092 50102 189750 50130
rect 190472 50102 190762 50130
rect 187516 47864 187568 47870
rect 187516 47806 187568 47812
rect 187332 3596 187384 3602
rect 187332 3538 187384 3544
rect 186148 3454 186452 3482
rect 186148 480 186176 3454
rect 187344 480 187372 3538
rect 187712 3534 187740 50102
rect 189092 3534 189120 50102
rect 187700 3528 187752 3534
rect 187700 3470 187752 3476
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 189080 3528 189132 3534
rect 189080 3470 189132 3476
rect 189724 3528 189776 3534
rect 189724 3470 189776 3476
rect 188540 480 188568 3470
rect 189736 480 189764 3470
rect 190472 490 190500 50102
rect 191852 16574 191880 50116
rect 192970 50102 193168 50130
rect 191852 16546 192064 16574
rect 190656 598 190868 626
rect 190656 490 190684 598
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 462 190684 490
rect 190840 480 190868 598
rect 192036 480 192064 16546
rect 193140 3074 193168 50102
rect 194060 47802 194088 50116
rect 194612 50102 195178 50130
rect 195992 50102 196282 50130
rect 193312 47796 193364 47802
rect 193312 47738 193364 47744
rect 194048 47796 194100 47802
rect 194048 47738 194100 47744
rect 193324 16574 193352 47738
rect 193324 16546 194456 16574
rect 193140 3046 193260 3074
rect 193232 480 193260 3046
rect 194428 480 194456 16546
rect 194612 3534 194640 50102
rect 194600 3528 194652 3534
rect 194600 3470 194652 3476
rect 195612 3528 195664 3534
rect 195612 3470 195664 3476
rect 195624 480 195652 3470
rect 195992 3466 196020 50102
rect 197372 16574 197400 50116
rect 198490 50102 198688 50130
rect 197372 16546 197952 16574
rect 195980 3460 196032 3466
rect 195980 3402 196032 3408
rect 196808 3460 196860 3466
rect 196808 3402 196860 3408
rect 196820 480 196848 3402
rect 197924 480 197952 16546
rect 198660 3534 198688 50102
rect 199580 46986 199608 50116
rect 200698 50102 201448 50130
rect 199568 46980 199620 46986
rect 199568 46922 199620 46928
rect 200212 46980 200264 46986
rect 200212 46922 200264 46928
rect 200224 16574 200252 46922
rect 200224 16546 200344 16574
rect 198648 3528 198700 3534
rect 198648 3470 198700 3476
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 199120 480 199148 3470
rect 200316 480 200344 16546
rect 201420 3482 201448 50102
rect 201512 50102 201802 50130
rect 201512 3602 201540 50102
rect 201500 3596 201552 3602
rect 201500 3538 201552 3544
rect 202696 3596 202748 3602
rect 202696 3538 202748 3544
rect 201420 3454 201540 3482
rect 201512 480 201540 3454
rect 202708 480 202736 3538
rect 202800 3534 202828 50116
rect 203918 50102 204208 50130
rect 205022 50102 205588 50130
rect 204180 47818 204208 50102
rect 204180 47790 204392 47818
rect 204364 16574 204392 47790
rect 204364 16546 205128 16574
rect 202788 3528 202840 3534
rect 202788 3470 202840 3476
rect 203892 3528 203944 3534
rect 203892 3470 203944 3476
rect 203904 480 203932 3470
rect 205100 480 205128 16546
rect 205560 3534 205588 50102
rect 206112 47870 206140 50116
rect 206100 47864 206152 47870
rect 206100 47806 206152 47812
rect 206928 47864 206980 47870
rect 206928 47806 206980 47812
rect 206940 3534 206968 47806
rect 207216 47326 207244 50116
rect 207204 47320 207256 47326
rect 207204 47262 207256 47268
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 206192 3528 206244 3534
rect 206192 3470 206244 3476
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 207388 3528 207440 3534
rect 207388 3470 207440 3476
rect 206204 480 206232 3470
rect 207400 480 207428 3470
rect 208320 3262 208348 50116
rect 209438 50102 209728 50130
rect 210542 50102 211108 50130
rect 208492 47320 208544 47326
rect 208492 47262 208544 47268
rect 208504 16574 208532 47262
rect 208504 16546 208624 16574
rect 208308 3256 208360 3262
rect 208308 3198 208360 3204
rect 208596 480 208624 16546
rect 209700 4146 209728 50102
rect 209688 4140 209740 4146
rect 209688 4082 209740 4088
rect 210976 4140 211028 4146
rect 210976 4082 211028 4088
rect 209780 3256 209832 3262
rect 209780 3198 209832 3204
rect 209792 480 209820 3198
rect 210988 480 211016 4082
rect 211080 3534 211108 50102
rect 211632 47802 211660 50116
rect 212736 47938 212764 50116
rect 212724 47932 212776 47938
rect 212724 47874 212776 47880
rect 211620 47796 211672 47802
rect 211620 47738 211672 47744
rect 212724 47796 212776 47802
rect 212724 47738 212776 47744
rect 212736 16574 212764 47738
rect 212736 16546 213408 16574
rect 211068 3528 211120 3534
rect 211068 3470 211120 3476
rect 212172 3528 212224 3534
rect 212172 3470 212224 3476
rect 212184 480 212212 3470
rect 213380 480 213408 16546
rect 213840 2990 213868 50116
rect 214866 50102 215248 50130
rect 215970 50102 216628 50130
rect 214012 47932 214064 47938
rect 214012 47874 214064 47880
rect 214024 16574 214052 47874
rect 214024 16546 214512 16574
rect 213828 2984 213880 2990
rect 213828 2926 213880 2932
rect 214484 480 214512 16546
rect 215220 3534 215248 50102
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 216600 3466 216628 50102
rect 217060 47870 217088 50116
rect 217048 47864 217100 47870
rect 217048 47806 217100 47812
rect 217968 47864 218020 47870
rect 217968 47806 218020 47812
rect 217980 3534 218008 47806
rect 218164 47666 218192 50116
rect 218152 47660 218204 47666
rect 218152 47602 218204 47608
rect 219268 46986 219296 50116
rect 220386 50102 220768 50130
rect 219348 47660 219400 47666
rect 219348 47602 219400 47608
rect 219256 46980 219308 46986
rect 219256 46922 219308 46928
rect 219360 3602 219388 47602
rect 220084 46980 220136 46986
rect 220084 46922 220136 46928
rect 219348 3596 219400 3602
rect 219348 3538 219400 3544
rect 220096 3534 220124 46922
rect 220452 3596 220504 3602
rect 220452 3538 220504 3544
rect 216864 3528 216916 3534
rect 216864 3470 216916 3476
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 219256 3528 219308 3534
rect 219256 3470 219308 3476
rect 220084 3528 220136 3534
rect 220084 3470 220136 3476
rect 216588 3460 216640 3466
rect 216588 3402 216640 3408
rect 215668 2984 215720 2990
rect 215668 2926 215720 2932
rect 215680 480 215708 2926
rect 216876 480 216904 3470
rect 218060 3460 218112 3466
rect 218060 3402 218112 3408
rect 218072 480 218100 3402
rect 219268 480 219296 3470
rect 220464 480 220492 3538
rect 220740 3330 220768 50102
rect 221476 47666 221504 50116
rect 222580 47870 222608 50116
rect 222568 47864 222620 47870
rect 222568 47806 222620 47812
rect 223488 47864 223540 47870
rect 223488 47806 223540 47812
rect 221464 47660 221516 47666
rect 221464 47602 221516 47608
rect 222844 47660 222896 47666
rect 222844 47602 222896 47608
rect 222856 3534 222884 47602
rect 223500 3602 223528 47806
rect 223684 47666 223712 50116
rect 224802 50102 224908 50130
rect 223672 47660 223724 47666
rect 223672 47602 223724 47608
rect 224776 47660 224828 47666
rect 224776 47602 224828 47608
rect 223488 3596 223540 3602
rect 223488 3538 223540 3544
rect 221556 3528 221608 3534
rect 221556 3470 221608 3476
rect 222844 3528 222896 3534
rect 222844 3470 222896 3476
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 220728 3324 220780 3330
rect 220728 3266 220780 3272
rect 221568 480 221596 3470
rect 222752 3324 222804 3330
rect 222752 3266 222804 3272
rect 222764 480 222792 3266
rect 223960 480 223988 3470
rect 224788 2990 224816 47602
rect 224880 3466 224908 50102
rect 225800 47802 225828 50116
rect 226904 47870 226932 50116
rect 228008 47870 228036 50116
rect 229112 47870 229140 50116
rect 230230 50102 230428 50130
rect 231334 50102 231808 50130
rect 226892 47864 226944 47870
rect 226892 47806 226944 47812
rect 227628 47864 227680 47870
rect 227628 47806 227680 47812
rect 227996 47864 228048 47870
rect 227996 47806 228048 47812
rect 229008 47864 229060 47870
rect 229008 47806 229060 47812
rect 229100 47864 229152 47870
rect 229100 47806 229152 47812
rect 225788 47796 225840 47802
rect 225788 47738 225840 47744
rect 225144 3596 225196 3602
rect 225144 3538 225196 3544
rect 224868 3460 224920 3466
rect 224868 3402 224920 3408
rect 224776 2984 224828 2990
rect 224776 2926 224828 2932
rect 225156 480 225184 3538
rect 227640 3534 227668 47806
rect 227812 47796 227864 47802
rect 227812 47738 227864 47744
rect 227824 16574 227852 47738
rect 227824 16546 228312 16574
rect 227628 3528 227680 3534
rect 227628 3470 227680 3476
rect 227536 3460 227588 3466
rect 227536 3402 227588 3408
rect 226340 2984 226392 2990
rect 226340 2926 226392 2932
rect 226352 480 226380 2926
rect 227548 480 227576 3402
rect 228284 490 228312 16546
rect 229020 4146 229048 47806
rect 229008 4140 229060 4146
rect 229008 4082 229060 4088
rect 229836 3528 229888 3534
rect 229836 3470 229888 3476
rect 228560 598 228772 626
rect 228560 490 228588 598
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 462 228588 490
rect 228744 480 228772 598
rect 229848 480 229876 3470
rect 230400 3194 230428 50102
rect 231032 4140 231084 4146
rect 231032 4082 231084 4088
rect 230388 3188 230440 3194
rect 230388 3130 230440 3136
rect 231044 480 231072 4082
rect 231780 3466 231808 50102
rect 232424 47870 232452 50116
rect 233528 47870 233556 50116
rect 234632 47870 234660 50116
rect 235750 50102 235948 50130
rect 236854 50102 237328 50130
rect 231952 47864 232004 47870
rect 231952 47806 232004 47812
rect 232412 47864 232464 47870
rect 232412 47806 232464 47812
rect 233148 47864 233200 47870
rect 233148 47806 233200 47812
rect 233516 47864 233568 47870
rect 233516 47806 233568 47812
rect 234528 47864 234580 47870
rect 234528 47806 234580 47812
rect 234620 47864 234672 47870
rect 234620 47806 234672 47812
rect 231964 16574 231992 47806
rect 231964 16546 232268 16574
rect 231768 3460 231820 3466
rect 231768 3402 231820 3408
rect 232240 480 232268 16546
rect 233160 3534 233188 47806
rect 233148 3528 233200 3534
rect 233148 3470 233200 3476
rect 234540 3194 234568 47806
rect 235920 3738 235948 50102
rect 237300 4146 237328 50102
rect 237852 47870 237880 50116
rect 237472 47864 237524 47870
rect 237472 47806 237524 47812
rect 237840 47864 237892 47870
rect 237840 47806 237892 47812
rect 238668 47864 238720 47870
rect 238668 47806 238720 47812
rect 237484 16574 237512 47806
rect 237484 16546 237696 16574
rect 237288 4140 237340 4146
rect 237288 4082 237340 4088
rect 235908 3732 235960 3738
rect 235908 3674 235960 3680
rect 235816 3528 235868 3534
rect 235816 3470 235868 3476
rect 234620 3460 234672 3466
rect 234620 3402 234672 3408
rect 233424 3188 233476 3194
rect 233424 3130 233476 3136
rect 234528 3188 234580 3194
rect 234528 3130 234580 3136
rect 233436 480 233464 3130
rect 234632 480 234660 3402
rect 235828 480 235856 3470
rect 237012 3188 237064 3194
rect 237012 3130 237064 3136
rect 237024 480 237052 3130
rect 237668 490 237696 16546
rect 238680 3670 238708 47806
rect 238956 47734 238984 50116
rect 240060 47870 240088 50116
rect 241178 50102 241468 50130
rect 242282 50102 242848 50130
rect 240048 47864 240100 47870
rect 240048 47806 240100 47812
rect 240784 47864 240836 47870
rect 240784 47806 240836 47812
rect 238944 47728 238996 47734
rect 238944 47670 238996 47676
rect 240048 47728 240100 47734
rect 240048 47670 240100 47676
rect 239312 3732 239364 3738
rect 239312 3674 239364 3680
rect 238668 3664 238720 3670
rect 238668 3606 238720 3612
rect 237944 598 238156 626
rect 237944 490 237972 598
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 237668 462 237972 490
rect 238128 480 238156 598
rect 239324 480 239352 3674
rect 240060 3194 240088 47670
rect 240508 4140 240560 4146
rect 240508 4082 240560 4088
rect 240048 3188 240100 3194
rect 240048 3130 240100 3136
rect 240520 480 240548 4082
rect 240796 3534 240824 47806
rect 240784 3528 240836 3534
rect 240784 3470 240836 3476
rect 241440 3466 241468 50102
rect 241704 3664 241756 3670
rect 241704 3606 241756 3612
rect 241428 3460 241480 3466
rect 241428 3402 241480 3408
rect 241716 480 241744 3606
rect 242820 3602 242848 50102
rect 243372 47802 243400 50116
rect 244476 47870 244504 50116
rect 245488 50102 245594 50130
rect 246698 50102 246988 50130
rect 247802 50102 248368 50130
rect 244464 47864 244516 47870
rect 244464 47806 244516 47812
rect 243360 47796 243412 47802
rect 243360 47738 243412 47744
rect 245488 4010 245516 50102
rect 245568 47864 245620 47870
rect 245568 47806 245620 47812
rect 245476 4004 245528 4010
rect 245476 3946 245528 3952
rect 242808 3596 242860 3602
rect 242808 3538 242860 3544
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 242900 3188 242952 3194
rect 242900 3130 242952 3136
rect 242912 480 242940 3130
rect 244108 480 244136 3470
rect 245200 3460 245252 3466
rect 245200 3402 245252 3408
rect 245212 480 245240 3402
rect 245580 3262 245608 47806
rect 246304 47796 246356 47802
rect 246304 47738 246356 47744
rect 245568 3256 245620 3262
rect 245568 3198 245620 3204
rect 246316 3194 246344 47738
rect 246396 3596 246448 3602
rect 246396 3538 246448 3544
rect 246304 3188 246356 3194
rect 246304 3130 246356 3136
rect 246408 480 246436 3538
rect 246960 3534 246988 50102
rect 248340 3874 248368 50102
rect 248892 47870 248920 50116
rect 249904 47870 249932 50116
rect 251022 50102 251128 50130
rect 252126 50102 252508 50130
rect 253230 50102 253888 50130
rect 248880 47864 248932 47870
rect 248880 47806 248932 47812
rect 249708 47864 249760 47870
rect 249708 47806 249760 47812
rect 249892 47864 249944 47870
rect 249892 47806 249944 47812
rect 250996 47864 251048 47870
rect 250996 47806 251048 47812
rect 248328 3868 248380 3874
rect 248328 3810 248380 3816
rect 246948 3528 247000 3534
rect 246948 3470 247000 3476
rect 249720 3466 249748 47806
rect 249984 4004 250036 4010
rect 249984 3946 250036 3952
rect 249708 3460 249760 3466
rect 249708 3402 249760 3408
rect 247592 3188 247644 3194
rect 247592 3130 247644 3136
rect 248788 3188 248840 3194
rect 248788 3130 248840 3136
rect 247604 480 247632 3130
rect 248800 480 248828 3130
rect 249996 480 250024 3946
rect 251008 3262 251036 47806
rect 251100 3602 251128 50102
rect 252376 3868 252428 3874
rect 252376 3810 252428 3816
rect 251088 3596 251140 3602
rect 251088 3538 251140 3544
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 250996 3256 251048 3262
rect 250996 3198 251048 3204
rect 251192 480 251220 3470
rect 252388 480 252416 3810
rect 252480 3330 252508 50102
rect 253860 4078 253888 50102
rect 254320 47870 254348 50116
rect 255424 47870 255452 50116
rect 256542 50102 256648 50130
rect 257646 50102 258028 50130
rect 258750 50102 259408 50130
rect 254308 47864 254360 47870
rect 254308 47806 254360 47812
rect 255228 47864 255280 47870
rect 255228 47806 255280 47812
rect 255412 47864 255464 47870
rect 255412 47806 255464 47812
rect 256516 47864 256568 47870
rect 256516 47806 256568 47812
rect 253848 4072 253900 4078
rect 253848 4014 253900 4020
rect 253480 3460 253532 3466
rect 253480 3402 253532 3408
rect 252468 3324 252520 3330
rect 252468 3266 252520 3272
rect 253492 480 253520 3402
rect 254676 3256 254728 3262
rect 254676 3198 254728 3204
rect 254688 480 254716 3198
rect 255240 2922 255268 47806
rect 256528 4146 256556 47806
rect 256516 4140 256568 4146
rect 256516 4082 256568 4088
rect 255872 3596 255924 3602
rect 255872 3538 255924 3544
rect 255228 2916 255280 2922
rect 255228 2858 255280 2864
rect 255884 480 255912 3538
rect 256620 3534 256648 50102
rect 258000 3670 258028 50102
rect 258264 4072 258316 4078
rect 258264 4014 258316 4020
rect 257988 3664 258040 3670
rect 257988 3606 258040 3612
rect 256608 3528 256660 3534
rect 256608 3470 256660 3476
rect 257068 3324 257120 3330
rect 257068 3266 257120 3272
rect 257080 480 257108 3266
rect 258276 480 258304 4014
rect 259380 3466 259408 50102
rect 259840 47598 259868 50116
rect 260944 47870 260972 50116
rect 261970 50102 262168 50130
rect 263074 50102 263548 50130
rect 264178 50102 264928 50130
rect 260932 47864 260984 47870
rect 260932 47806 260984 47812
rect 259828 47592 259880 47598
rect 259828 47534 259880 47540
rect 260748 47592 260800 47598
rect 260748 47534 260800 47540
rect 260656 4140 260708 4146
rect 260656 4082 260708 4088
rect 259368 3460 259420 3466
rect 259368 3402 259420 3408
rect 259460 2916 259512 2922
rect 259460 2858 259512 2864
rect 259472 480 259500 2858
rect 260668 480 260696 4082
rect 260760 3330 260788 47534
rect 262140 4146 262168 50102
rect 262128 4140 262180 4146
rect 262128 4082 262180 4088
rect 262956 3664 263008 3670
rect 262956 3606 263008 3612
rect 261760 3528 261812 3534
rect 261760 3470 261812 3476
rect 260748 3324 260800 3330
rect 260748 3266 260800 3272
rect 261772 480 261800 3470
rect 262968 480 262996 3606
rect 263520 3058 263548 50102
rect 264244 47864 264296 47870
rect 264244 47806 264296 47812
rect 264152 3460 264204 3466
rect 264152 3402 264204 3408
rect 263508 3052 263560 3058
rect 263508 2994 263560 3000
rect 264164 480 264192 3402
rect 264256 3194 264284 47806
rect 264900 4010 264928 50102
rect 265268 47598 265296 50116
rect 266372 47666 266400 50116
rect 267490 50102 267596 50130
rect 268594 50102 269068 50130
rect 269698 50102 270448 50130
rect 266360 47660 266412 47666
rect 266360 47602 266412 47608
rect 265256 47592 265308 47598
rect 265256 47534 265308 47540
rect 264888 4004 264940 4010
rect 264888 3946 264940 3952
rect 267568 3466 267596 50102
rect 267648 47660 267700 47666
rect 267648 47602 267700 47608
rect 267660 3738 267688 47602
rect 267740 4140 267792 4146
rect 267740 4082 267792 4088
rect 267648 3732 267700 3738
rect 267648 3674 267700 3680
rect 267556 3460 267608 3466
rect 267556 3402 267608 3408
rect 265348 3324 265400 3330
rect 265348 3266 265400 3272
rect 264244 3188 264296 3194
rect 264244 3130 264296 3136
rect 265360 480 265388 3266
rect 266544 3188 266596 3194
rect 266544 3130 266596 3136
rect 266556 480 266584 3130
rect 267752 480 267780 4082
rect 269040 3534 269068 50102
rect 270040 4004 270092 4010
rect 270040 3946 270092 3952
rect 269028 3528 269080 3534
rect 269028 3470 269080 3476
rect 268844 3052 268896 3058
rect 268844 2994 268896 3000
rect 268856 480 268884 2994
rect 270052 480 270080 3946
rect 270420 2990 270448 50102
rect 270788 47870 270816 50116
rect 270776 47864 270828 47870
rect 270776 47806 270828 47812
rect 271788 47864 271840 47870
rect 271788 47806 271840 47812
rect 270592 47592 270644 47598
rect 270592 47534 270644 47540
rect 270604 16574 270632 47534
rect 270604 16546 270816 16574
rect 270408 2984 270460 2990
rect 270408 2926 270460 2932
rect 270788 490 270816 16546
rect 271800 3330 271828 47806
rect 271892 47054 271920 50116
rect 272918 50102 273208 50130
rect 274022 50102 274588 50130
rect 271880 47048 271932 47054
rect 271880 46990 271932 46996
rect 272432 3732 272484 3738
rect 272432 3674 272484 3680
rect 271788 3324 271840 3330
rect 271788 3266 271840 3272
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 3674
rect 273180 3194 273208 50102
rect 274560 3874 274588 50102
rect 275112 47598 275140 50116
rect 276216 47666 276244 50116
rect 277228 50102 277334 50130
rect 278438 50102 278728 50130
rect 279542 50102 280108 50130
rect 276204 47660 276256 47666
rect 276204 47602 276256 47608
rect 275100 47592 275152 47598
rect 275100 47534 275152 47540
rect 275928 47592 275980 47598
rect 275928 47534 275980 47540
rect 274548 3868 274600 3874
rect 274548 3810 274600 3816
rect 275940 3738 275968 47534
rect 275928 3732 275980 3738
rect 275928 3674 275980 3680
rect 274824 3528 274876 3534
rect 274824 3470 274876 3476
rect 273628 3460 273680 3466
rect 273628 3402 273680 3408
rect 273168 3188 273220 3194
rect 273168 3130 273220 3136
rect 273640 480 273668 3402
rect 274836 480 274864 3470
rect 277228 3466 277256 50102
rect 277308 47660 277360 47666
rect 277308 47602 277360 47608
rect 277320 3670 277348 47602
rect 277492 47048 277544 47054
rect 277492 46990 277544 46996
rect 277504 16574 277532 46990
rect 277504 16546 278360 16574
rect 277308 3664 277360 3670
rect 277308 3606 277360 3612
rect 277216 3460 277268 3466
rect 277216 3402 277268 3408
rect 277124 3324 277176 3330
rect 277124 3266 277176 3272
rect 276020 2984 276072 2990
rect 276020 2926 276072 2932
rect 276032 480 276060 2926
rect 277136 480 277164 3266
rect 278332 480 278360 16546
rect 278700 3330 278728 50102
rect 278688 3324 278740 3330
rect 278688 3266 278740 3272
rect 279516 3188 279568 3194
rect 279516 3130 279568 3136
rect 279528 480 279556 3130
rect 280080 2990 280108 50102
rect 280632 47598 280660 50116
rect 281736 47870 281764 50116
rect 281724 47864 281776 47870
rect 281724 47806 281776 47812
rect 282736 47864 282788 47870
rect 282736 47806 282788 47812
rect 280620 47592 280672 47598
rect 280620 47534 280672 47540
rect 281448 47592 281500 47598
rect 281448 47534 281500 47540
rect 281460 4010 281488 47534
rect 282748 4146 282776 47806
rect 282736 4140 282788 4146
rect 282736 4082 282788 4088
rect 281448 4004 281500 4010
rect 281448 3946 281500 3952
rect 280712 3868 280764 3874
rect 280712 3810 280764 3816
rect 280068 2984 280120 2990
rect 280068 2926 280120 2932
rect 280724 480 280752 3810
rect 281908 3732 281960 3738
rect 281908 3674 281960 3680
rect 281920 480 281948 3674
rect 282840 3602 282868 50116
rect 283958 50102 284248 50130
rect 284970 50102 285628 50130
rect 284220 3738 284248 50102
rect 284208 3732 284260 3738
rect 284208 3674 284260 3680
rect 285600 3670 285628 50102
rect 286060 47870 286088 50116
rect 287164 47870 287192 50116
rect 286048 47864 286100 47870
rect 286048 47806 286100 47812
rect 286968 47864 287020 47870
rect 286968 47806 287020 47812
rect 287152 47864 287204 47870
rect 287152 47806 287204 47812
rect 286980 3806 287008 47806
rect 287796 4004 287848 4010
rect 287796 3946 287848 3952
rect 286968 3800 287020 3806
rect 286968 3742 287020 3748
rect 283104 3664 283156 3670
rect 283104 3606 283156 3612
rect 285588 3664 285640 3670
rect 285588 3606 285640 3612
rect 282828 3596 282880 3602
rect 282828 3538 282880 3544
rect 283116 480 283144 3606
rect 284300 3460 284352 3466
rect 284300 3402 284352 3408
rect 284312 480 284340 3402
rect 285404 3324 285456 3330
rect 285404 3266 285456 3272
rect 285416 480 285444 3266
rect 286600 2984 286652 2990
rect 286600 2926 286652 2932
rect 286612 480 286640 2926
rect 287808 480 287836 3946
rect 288268 3330 288296 50116
rect 289386 50102 289768 50130
rect 290490 50102 291148 50130
rect 288348 47864 288400 47870
rect 288348 47806 288400 47812
rect 288256 3324 288308 3330
rect 288256 3266 288308 3272
rect 288360 2922 288388 47806
rect 288992 4140 289044 4146
rect 288992 4082 289044 4088
rect 288348 2916 288400 2922
rect 288348 2858 288400 2864
rect 289004 480 289032 4082
rect 289740 3534 289768 50102
rect 290188 3596 290240 3602
rect 290188 3538 290240 3544
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 290200 480 290228 3538
rect 291120 3058 291148 50102
rect 291580 47870 291608 50116
rect 292684 47870 292712 50116
rect 293802 50102 293908 50130
rect 294906 50102 295288 50130
rect 296010 50102 296668 50130
rect 291568 47864 291620 47870
rect 291568 47806 291620 47812
rect 292488 47864 292540 47870
rect 292488 47806 292540 47812
rect 292672 47864 292724 47870
rect 292672 47806 292724 47812
rect 293776 47864 293828 47870
rect 293776 47806 293828 47812
rect 292500 3874 292528 47806
rect 293788 4010 293816 47806
rect 293776 4004 293828 4010
rect 293776 3946 293828 3952
rect 292488 3868 292540 3874
rect 292488 3810 292540 3816
rect 293684 3800 293736 3806
rect 293684 3742 293736 3748
rect 291384 3732 291436 3738
rect 291384 3674 291436 3680
rect 291108 3052 291160 3058
rect 291108 2994 291160 3000
rect 291396 480 291424 3674
rect 292580 3664 292632 3670
rect 292580 3606 292632 3612
rect 292592 480 292620 3606
rect 293696 480 293724 3742
rect 293880 3670 293908 50102
rect 295260 3738 295288 50102
rect 295248 3732 295300 3738
rect 295248 3674 295300 3680
rect 293868 3664 293920 3670
rect 293868 3606 293920 3612
rect 296640 3466 296668 50102
rect 297008 47870 297036 50116
rect 296996 47864 297048 47870
rect 296996 47806 297048 47812
rect 298008 47864 298060 47870
rect 298008 47806 298060 47812
rect 297272 3528 297324 3534
rect 297272 3470 297324 3476
rect 296628 3460 296680 3466
rect 296628 3402 296680 3408
rect 296076 3324 296128 3330
rect 296076 3266 296128 3272
rect 294880 2916 294932 2922
rect 294880 2858 294932 2864
rect 294892 480 294920 2858
rect 296088 480 296116 3266
rect 297284 480 297312 3470
rect 298020 3330 298048 47806
rect 298112 47326 298140 50116
rect 299230 50102 299428 50130
rect 300334 50102 300808 50130
rect 298100 47320 298152 47326
rect 298100 47262 298152 47268
rect 299296 47320 299348 47326
rect 299296 47262 299348 47268
rect 299308 3534 299336 47262
rect 299400 3602 299428 50102
rect 300780 6914 300808 50102
rect 301424 47870 301452 50116
rect 302528 47870 302556 50116
rect 303632 47870 303660 50116
rect 304750 50102 304856 50130
rect 305854 50102 306328 50130
rect 301412 47864 301464 47870
rect 301412 47806 301464 47812
rect 302148 47864 302200 47870
rect 302148 47806 302200 47812
rect 302516 47864 302568 47870
rect 302516 47806 302568 47812
rect 303528 47864 303580 47870
rect 303528 47806 303580 47812
rect 303620 47864 303672 47870
rect 303620 47806 303672 47812
rect 300688 6886 300808 6914
rect 299664 3868 299716 3874
rect 299664 3810 299716 3816
rect 299388 3596 299440 3602
rect 299388 3538 299440 3544
rect 299296 3528 299348 3534
rect 299296 3470 299348 3476
rect 298008 3324 298060 3330
rect 298008 3266 298060 3272
rect 298468 3052 298520 3058
rect 298468 2994 298520 3000
rect 298480 480 298508 2994
rect 299676 480 299704 3810
rect 300688 3398 300716 6886
rect 300768 4004 300820 4010
rect 300768 3946 300820 3952
rect 300676 3392 300728 3398
rect 300676 3334 300728 3340
rect 300780 480 300808 3946
rect 302160 3670 302188 47806
rect 303540 3942 303568 47806
rect 303528 3936 303580 3942
rect 303528 3878 303580 3884
rect 303160 3732 303212 3738
rect 303160 3674 303212 3680
rect 301964 3664 302016 3670
rect 301964 3606 302016 3612
rect 302148 3664 302200 3670
rect 302148 3606 302200 3612
rect 301976 480 302004 3606
rect 303172 480 303200 3674
rect 304828 3466 304856 50102
rect 304908 47864 304960 47870
rect 304908 47806 304960 47812
rect 304920 4078 304948 47806
rect 304908 4072 304960 4078
rect 304908 4014 304960 4020
rect 306300 3738 306328 50102
rect 306944 47802 306972 50116
rect 307956 47870 307984 50116
rect 307944 47864 307996 47870
rect 307944 47806 307996 47812
rect 308956 47864 309008 47870
rect 308956 47806 309008 47812
rect 306932 47796 306984 47802
rect 306932 47738 306984 47744
rect 307668 47796 307720 47802
rect 307668 47738 307720 47744
rect 306288 3732 306340 3738
rect 306288 3674 306340 3680
rect 307680 3534 307708 47738
rect 308968 3874 308996 47806
rect 308956 3868 309008 3874
rect 308956 3810 309008 3816
rect 309060 3806 309088 50116
rect 310178 50102 310468 50130
rect 311282 50102 311848 50130
rect 309048 3800 309100 3806
rect 309048 3742 309100 3748
rect 310244 3664 310296 3670
rect 310244 3606 310296 3612
rect 307944 3596 307996 3602
rect 307944 3538 307996 3544
rect 306748 3528 306800 3534
rect 306748 3470 306800 3476
rect 307668 3528 307720 3534
rect 307668 3470 307720 3476
rect 304356 3460 304408 3466
rect 304356 3402 304408 3408
rect 304816 3460 304868 3466
rect 304816 3402 304868 3408
rect 304368 480 304396 3402
rect 305552 3324 305604 3330
rect 305552 3266 305604 3272
rect 305564 480 305592 3266
rect 306760 480 306788 3470
rect 307956 480 307984 3538
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 310256 480 310284 3606
rect 310440 3602 310468 50102
rect 311820 4010 311848 50102
rect 312372 47870 312400 50116
rect 312360 47864 312412 47870
rect 312360 47806 312412 47812
rect 313188 47864 313240 47870
rect 313188 47806 313240 47812
rect 312636 4072 312688 4078
rect 312636 4014 312688 4020
rect 311808 4004 311860 4010
rect 311808 3946 311860 3952
rect 311440 3936 311492 3942
rect 311440 3878 311492 3884
rect 310428 3596 310480 3602
rect 310428 3538 310480 3544
rect 311452 480 311480 3878
rect 312648 480 312676 4014
rect 313200 3670 313228 47806
rect 313476 47666 313504 50116
rect 314488 50102 314594 50130
rect 315698 50102 315988 50130
rect 316802 50102 317368 50130
rect 313464 47660 313516 47666
rect 313464 47602 313516 47608
rect 313188 3664 313240 3670
rect 313188 3606 313240 3612
rect 314488 3466 314516 50102
rect 314568 47660 314620 47666
rect 314568 47602 314620 47608
rect 314580 4078 314608 47602
rect 314568 4072 314620 4078
rect 314568 4014 314620 4020
rect 315960 3738 315988 50102
rect 317340 4010 317368 50102
rect 317892 47870 317920 50116
rect 317880 47864 317932 47870
rect 317880 47806 317932 47812
rect 318708 47864 318760 47870
rect 318708 47806 318760 47812
rect 317328 4004 317380 4010
rect 317328 3946 317380 3952
rect 318720 3874 318748 47806
rect 318996 47802 319024 50116
rect 318984 47796 319036 47802
rect 318984 47738 319036 47744
rect 317328 3868 317380 3874
rect 317328 3810 317380 3816
rect 318708 3868 318760 3874
rect 318708 3810 318760 3816
rect 315028 3732 315080 3738
rect 315028 3674 315080 3680
rect 315948 3732 316000 3738
rect 315948 3674 316000 3680
rect 313832 3460 313884 3466
rect 313832 3402 313884 3408
rect 314476 3460 314528 3466
rect 314476 3402 314528 3408
rect 313844 480 313872 3402
rect 315040 480 315068 3674
rect 316224 3528 316276 3534
rect 316224 3470 316276 3476
rect 316236 480 316264 3470
rect 317340 480 317368 3810
rect 318524 3800 318576 3806
rect 318524 3742 318576 3748
rect 318536 480 318564 3742
rect 319720 3596 319772 3602
rect 319720 3538 319772 3544
rect 319732 480 319760 3538
rect 320008 3398 320036 50116
rect 321126 50102 321508 50130
rect 322230 50102 322888 50130
rect 320088 47796 320140 47802
rect 320088 47738 320140 47744
rect 320100 3806 320128 47738
rect 320916 4072 320968 4078
rect 320916 4014 320968 4020
rect 320088 3800 320140 3806
rect 320088 3742 320140 3748
rect 319996 3392 320048 3398
rect 319996 3334 320048 3340
rect 320928 480 320956 4014
rect 321480 3534 321508 50102
rect 322112 3664 322164 3670
rect 322112 3606 322164 3612
rect 321468 3528 321520 3534
rect 321468 3470 321520 3476
rect 322124 480 322152 3606
rect 322860 3602 322888 50102
rect 323320 47598 323348 50116
rect 324424 47870 324452 50116
rect 325542 50102 325648 50130
rect 326646 50102 327028 50130
rect 327750 50102 328408 50130
rect 324412 47864 324464 47870
rect 324412 47806 324464 47812
rect 325516 47864 325568 47870
rect 325516 47806 325568 47812
rect 323308 47592 323360 47598
rect 323308 47534 323360 47540
rect 324228 47592 324280 47598
rect 324228 47534 324280 47540
rect 324240 4146 324268 47534
rect 323308 4140 323360 4146
rect 323308 4082 323360 4088
rect 324228 4140 324280 4146
rect 324228 4082 324280 4088
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 323320 480 323348 4082
rect 325528 3738 325556 47806
rect 325620 3754 325648 50102
rect 327000 3942 327028 50102
rect 326804 3936 326856 3942
rect 326804 3878 326856 3884
rect 326988 3936 327040 3942
rect 326988 3878 327040 3884
rect 325516 3732 325568 3738
rect 325620 3726 325740 3754
rect 325516 3674 325568 3680
rect 325608 3664 325660 3670
rect 325608 3606 325660 3612
rect 324412 3460 324464 3466
rect 324412 3402 324464 3408
rect 324424 480 324452 3402
rect 325620 480 325648 3606
rect 325712 3466 325740 3726
rect 325700 3460 325752 3466
rect 325700 3402 325752 3408
rect 326816 480 326844 3878
rect 328380 3874 328408 50102
rect 328840 47870 328868 50116
rect 329944 47870 329972 50116
rect 328828 47864 328880 47870
rect 328828 47806 328880 47812
rect 329748 47864 329800 47870
rect 329748 47806 329800 47812
rect 329932 47864 329984 47870
rect 329932 47806 329984 47812
rect 328000 3868 328052 3874
rect 328000 3810 328052 3816
rect 328368 3868 328420 3874
rect 328368 3810 328420 3816
rect 328012 480 328040 3810
rect 329760 3806 329788 47806
rect 329196 3800 329248 3806
rect 329196 3742 329248 3748
rect 329748 3800 329800 3806
rect 329748 3742 329800 3748
rect 329208 480 329236 3742
rect 331048 3670 331076 50116
rect 332074 50102 332548 50130
rect 333178 50102 333928 50130
rect 331128 47864 331180 47870
rect 331128 47806 331180 47812
rect 331140 4078 331168 47806
rect 331128 4072 331180 4078
rect 331128 4014 331180 4020
rect 332520 4010 332548 50102
rect 333900 6914 333928 50102
rect 334268 47870 334296 50116
rect 335372 47870 335400 50116
rect 336490 50102 336596 50130
rect 337594 50102 338068 50130
rect 338698 50102 339448 50130
rect 334256 47864 334308 47870
rect 334256 47806 334308 47812
rect 335268 47864 335320 47870
rect 335268 47806 335320 47812
rect 335360 47864 335412 47870
rect 335360 47806 335412 47812
rect 333808 6886 333928 6914
rect 332508 4004 332560 4010
rect 332508 3946 332560 3952
rect 331036 3664 331088 3670
rect 331036 3606 331088 3612
rect 332692 3596 332744 3602
rect 332692 3538 332744 3544
rect 331588 3528 331640 3534
rect 331588 3470 331640 3476
rect 330392 3392 330444 3398
rect 330392 3334 330444 3340
rect 330404 480 330432 3334
rect 331600 480 331628 3470
rect 332704 480 332732 3538
rect 333808 3398 333836 6886
rect 333888 4140 333940 4146
rect 333888 4082 333940 4088
rect 333796 3392 333848 3398
rect 333796 3334 333848 3340
rect 333900 480 333928 4082
rect 335084 3732 335136 3738
rect 335084 3674 335136 3680
rect 335096 480 335124 3674
rect 335280 3670 335308 47806
rect 335268 3664 335320 3670
rect 335268 3606 335320 3612
rect 336568 3466 336596 50102
rect 336648 47864 336700 47870
rect 336648 47806 336700 47812
rect 336660 3738 336688 47806
rect 337476 3936 337528 3942
rect 337476 3878 337528 3884
rect 336648 3732 336700 3738
rect 336648 3674 336700 3680
rect 336280 3460 336332 3466
rect 336280 3402 336332 3408
rect 336556 3460 336608 3466
rect 336556 3402 336608 3408
rect 336292 480 336320 3402
rect 337488 480 337516 3878
rect 338040 3602 338068 50102
rect 339420 3874 339448 50102
rect 339788 47870 339816 50116
rect 339776 47864 339828 47870
rect 339776 47806 339828 47812
rect 340788 47864 340840 47870
rect 340788 47806 340840 47812
rect 338672 3868 338724 3874
rect 338672 3810 338724 3816
rect 339408 3868 339460 3874
rect 339408 3810 339460 3816
rect 338028 3596 338080 3602
rect 338028 3538 338080 3544
rect 338684 480 338712 3810
rect 339868 3800 339920 3806
rect 339868 3742 339920 3748
rect 339880 480 339908 3742
rect 340800 3262 340828 47806
rect 340892 47734 340920 50116
rect 342010 50102 342208 50130
rect 343114 50102 343588 50130
rect 340880 47728 340932 47734
rect 340880 47670 340932 47676
rect 342076 47728 342128 47734
rect 342076 47670 342128 47676
rect 342088 4078 342116 47670
rect 340972 4072 341024 4078
rect 340972 4014 341024 4020
rect 342076 4072 342128 4078
rect 342076 4014 342128 4020
rect 340788 3256 340840 3262
rect 340788 3198 340840 3204
rect 340984 480 341012 4014
rect 342180 3942 342208 50102
rect 343560 4146 343588 50102
rect 344112 47598 344140 50116
rect 344100 47592 344152 47598
rect 344100 47534 344152 47540
rect 344928 47592 344980 47598
rect 344928 47534 344980 47540
rect 343548 4140 343600 4146
rect 343548 4082 343600 4088
rect 343364 4004 343416 4010
rect 343364 3946 343416 3952
rect 342168 3936 342220 3942
rect 342168 3878 342220 3884
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 342180 480 342208 3470
rect 343376 480 343404 3946
rect 344940 3534 344968 47534
rect 345216 47462 345244 50116
rect 346228 50102 346334 50130
rect 347438 50102 347728 50130
rect 348542 50102 349108 50130
rect 345204 47456 345256 47462
rect 345204 47398 345256 47404
rect 346228 3670 346256 50102
rect 346308 47456 346360 47462
rect 346308 47398 346360 47404
rect 346320 4010 346348 47398
rect 346308 4004 346360 4010
rect 346308 3946 346360 3952
rect 347700 3806 347728 50102
rect 347688 3800 347740 3806
rect 347688 3742 347740 3748
rect 349080 3738 349108 50102
rect 349632 47598 349660 50116
rect 350736 47870 350764 50116
rect 350724 47864 350776 47870
rect 350724 47806 350776 47812
rect 351736 47864 351788 47870
rect 351736 47806 351788 47812
rect 349620 47592 349672 47598
rect 349620 47534 349672 47540
rect 350448 47592 350500 47598
rect 350448 47534 350500 47540
rect 350460 6914 350488 47534
rect 350368 6886 350488 6914
rect 346952 3732 347004 3738
rect 346952 3674 347004 3680
rect 349068 3732 349120 3738
rect 349068 3674 349120 3680
rect 345756 3664 345808 3670
rect 345756 3606 345808 3612
rect 346216 3664 346268 3670
rect 346216 3606 346268 3612
rect 344928 3528 344980 3534
rect 344928 3470 344980 3476
rect 344560 3392 344612 3398
rect 344560 3334 344612 3340
rect 344572 480 344600 3334
rect 345768 480 345796 3606
rect 346964 480 346992 3674
rect 349252 3596 349304 3602
rect 349252 3538 349304 3544
rect 348056 3460 348108 3466
rect 348056 3402 348108 3408
rect 348068 480 348096 3402
rect 349264 480 349292 3538
rect 350368 3330 350396 6886
rect 351748 3874 351776 47806
rect 350448 3868 350500 3874
rect 350448 3810 350500 3816
rect 351736 3868 351788 3874
rect 351736 3810 351788 3816
rect 350356 3324 350408 3330
rect 350356 3266 350408 3272
rect 350460 480 350488 3810
rect 351840 3466 351868 50116
rect 352958 50102 353248 50130
rect 354062 50102 354628 50130
rect 352840 4072 352892 4078
rect 352840 4014 352892 4020
rect 351828 3460 351880 3466
rect 351828 3402 351880 3408
rect 351644 3256 351696 3262
rect 351644 3198 351696 3204
rect 351656 480 351684 3198
rect 352852 480 352880 4014
rect 353220 3602 353248 50102
rect 354600 4078 354628 50102
rect 355060 47870 355088 50116
rect 355048 47864 355100 47870
rect 355048 47806 355100 47812
rect 355968 47864 356020 47870
rect 355968 47806 356020 47812
rect 355980 4146 356008 47806
rect 356164 47666 356192 50116
rect 356152 47660 356204 47666
rect 356152 47602 356204 47608
rect 355232 4140 355284 4146
rect 355232 4082 355284 4088
rect 355968 4140 356020 4146
rect 355968 4082 356020 4088
rect 354588 4072 354640 4078
rect 354588 4014 354640 4020
rect 354036 3936 354088 3942
rect 354036 3878 354088 3884
rect 353208 3596 353260 3602
rect 353208 3538 353260 3544
rect 354048 480 354076 3878
rect 355244 480 355272 4082
rect 356336 3528 356388 3534
rect 356336 3470 356388 3476
rect 356348 480 356376 3470
rect 357268 3398 357296 50116
rect 358386 50102 358768 50130
rect 359490 50102 360148 50130
rect 357348 47660 357400 47666
rect 357348 47602 357400 47608
rect 357256 3392 357308 3398
rect 357256 3334 357308 3340
rect 357360 3262 357388 47602
rect 357532 4004 357584 4010
rect 357532 3946 357584 3952
rect 357348 3256 357400 3262
rect 357348 3198 357400 3204
rect 357544 480 357572 3946
rect 358740 3806 358768 50102
rect 360120 3942 360148 50102
rect 360580 47870 360608 50116
rect 360568 47864 360620 47870
rect 360568 47806 360620 47812
rect 361488 47864 361540 47870
rect 361488 47806 361540 47812
rect 360108 3936 360160 3942
rect 360108 3878 360160 3884
rect 359924 3868 359976 3874
rect 359924 3810 359976 3816
rect 358728 3800 358780 3806
rect 358728 3742 358780 3748
rect 358728 3664 358780 3670
rect 358728 3606 358780 3612
rect 358740 480 358768 3606
rect 359936 480 359964 3810
rect 361500 3806 361528 47806
rect 361684 47666 361712 50116
rect 361672 47660 361724 47666
rect 361672 47602 361724 47608
rect 361488 3800 361540 3806
rect 361488 3742 361540 3748
rect 362788 3738 362816 50116
rect 363906 50102 364288 50130
rect 365010 50102 365668 50130
rect 362868 47660 362920 47666
rect 362868 47602 362920 47608
rect 362776 3732 362828 3738
rect 362776 3674 362828 3680
rect 361120 3528 361172 3534
rect 361120 3470 361172 3476
rect 361132 480 361160 3470
rect 362316 3324 362368 3330
rect 362316 3266 362368 3272
rect 362328 480 362356 3266
rect 362880 3262 362908 47602
rect 363512 3868 363564 3874
rect 363512 3810 363564 3816
rect 362868 3256 362920 3262
rect 362868 3198 362920 3204
rect 363524 480 363552 3810
rect 364260 3330 364288 50102
rect 365640 4010 365668 50102
rect 366100 47870 366128 50116
rect 367112 47870 367140 50116
rect 368230 50102 368428 50130
rect 369334 50102 369808 50130
rect 366088 47864 366140 47870
rect 366088 47806 366140 47812
rect 367008 47864 367060 47870
rect 367008 47806 367060 47812
rect 367100 47864 367152 47870
rect 367100 47806 367152 47812
rect 368296 47864 368348 47870
rect 368296 47806 368348 47812
rect 366916 4072 366968 4078
rect 366916 4014 366968 4020
rect 365628 4004 365680 4010
rect 365628 3946 365680 3952
rect 365812 3596 365864 3602
rect 365812 3538 365864 3544
rect 364616 3460 364668 3466
rect 364616 3402 364668 3408
rect 364248 3324 364300 3330
rect 364248 3266 364300 3272
rect 364628 480 364656 3402
rect 365824 480 365852 3538
rect 366928 1034 366956 4014
rect 367020 3874 367048 47806
rect 368204 4140 368256 4146
rect 368204 4082 368256 4088
rect 367008 3868 367060 3874
rect 367008 3810 367060 3816
rect 366928 1006 367048 1034
rect 367020 480 367048 1006
rect 368216 480 368244 4082
rect 368308 3602 368336 47806
rect 368296 3596 368348 3602
rect 368296 3538 368348 3544
rect 368400 3466 368428 50102
rect 368388 3460 368440 3466
rect 368388 3402 368440 3408
rect 369400 3392 369452 3398
rect 369400 3334 369452 3340
rect 369412 480 369440 3334
rect 369780 3194 369808 50102
rect 370424 47802 370452 50116
rect 371528 47870 371556 50116
rect 372632 47870 372660 50116
rect 373750 50102 373948 50130
rect 374854 50102 375328 50130
rect 371516 47864 371568 47870
rect 371516 47806 371568 47812
rect 372528 47864 372580 47870
rect 372528 47806 372580 47812
rect 372620 47864 372672 47870
rect 372620 47806 372672 47812
rect 373816 47864 373868 47870
rect 373816 47806 373868 47812
rect 370412 47796 370464 47802
rect 370412 47738 370464 47744
rect 371148 47796 371200 47802
rect 371148 47738 371200 47744
rect 371160 4146 371188 47738
rect 371148 4140 371200 4146
rect 371148 4082 371200 4088
rect 371700 3664 371752 3670
rect 371700 3606 371752 3612
rect 370596 3528 370648 3534
rect 370596 3470 370648 3476
rect 369768 3188 369820 3194
rect 369768 3130 369820 3136
rect 370608 480 370636 3470
rect 371712 480 371740 3606
rect 372540 3398 372568 47806
rect 373828 4078 373856 47806
rect 373816 4072 373868 4078
rect 373816 4014 373868 4020
rect 373920 3942 373948 50102
rect 372896 3936 372948 3942
rect 372896 3878 372948 3884
rect 373908 3936 373960 3942
rect 373908 3878 373960 3884
rect 372528 3392 372580 3398
rect 372528 3334 372580 3340
rect 372908 480 372936 3878
rect 374092 3800 374144 3806
rect 374092 3742 374144 3748
rect 374104 480 374132 3742
rect 375300 3670 375328 50102
rect 375944 47870 375972 50116
rect 377048 47870 377076 50116
rect 378152 47870 378180 50116
rect 379178 50102 379376 50130
rect 380282 50102 380848 50130
rect 375932 47864 375984 47870
rect 375932 47806 375984 47812
rect 376668 47864 376720 47870
rect 376668 47806 376720 47812
rect 377036 47864 377088 47870
rect 377036 47806 377088 47812
rect 378048 47864 378100 47870
rect 378048 47806 378100 47812
rect 378140 47864 378192 47870
rect 378140 47806 378192 47812
rect 376680 3738 376708 47806
rect 376484 3732 376536 3738
rect 376484 3674 376536 3680
rect 376668 3732 376720 3738
rect 376668 3674 376720 3680
rect 375288 3664 375340 3670
rect 375288 3606 375340 3612
rect 375288 3256 375340 3262
rect 375288 3198 375340 3204
rect 375300 480 375328 3198
rect 376496 480 376524 3674
rect 377680 3324 377732 3330
rect 377680 3266 377732 3272
rect 377692 480 377720 3266
rect 378060 3126 378088 47806
rect 378876 4004 378928 4010
rect 378876 3946 378928 3952
rect 378048 3120 378100 3126
rect 378048 3062 378100 3068
rect 378888 480 378916 3946
rect 379348 3534 379376 50102
rect 379428 47864 379480 47870
rect 379428 47806 379480 47812
rect 379336 3528 379388 3534
rect 379336 3470 379388 3476
rect 379440 3262 379468 47806
rect 379980 3868 380032 3874
rect 379980 3810 380032 3816
rect 379428 3256 379480 3262
rect 379428 3198 379480 3204
rect 379992 480 380020 3810
rect 380820 3806 380848 50102
rect 381372 47598 381400 50116
rect 382476 47870 382504 50116
rect 382464 47864 382516 47870
rect 382464 47806 382516 47812
rect 383476 47864 383528 47870
rect 383476 47806 383528 47812
rect 381360 47592 381412 47598
rect 381360 47534 381412 47540
rect 382188 47592 382240 47598
rect 382188 47534 382240 47540
rect 382200 4010 382228 47534
rect 382188 4004 382240 4010
rect 382188 3946 382240 3952
rect 383488 3874 383516 47806
rect 383476 3868 383528 3874
rect 383476 3810 383528 3816
rect 380808 3800 380860 3806
rect 380808 3742 380860 3748
rect 383580 3602 383608 50116
rect 384698 50102 384988 50130
rect 385802 50102 386368 50130
rect 384960 4146 384988 50102
rect 384764 4140 384816 4146
rect 384764 4082 384816 4088
rect 384948 4140 385000 4146
rect 384948 4082 385000 4088
rect 381176 3596 381228 3602
rect 381176 3538 381228 3544
rect 383568 3596 383620 3602
rect 383568 3538 383620 3544
rect 381188 480 381216 3538
rect 382372 3460 382424 3466
rect 382372 3402 382424 3408
rect 382384 480 382412 3402
rect 383568 3188 383620 3194
rect 383568 3130 383620 3136
rect 383580 480 383608 3130
rect 384776 480 384804 4082
rect 386340 3398 386368 50102
rect 386892 47870 386920 50116
rect 387996 47870 388024 50116
rect 389008 50102 389114 50130
rect 390126 50102 390508 50130
rect 391230 50102 391888 50130
rect 386880 47864 386932 47870
rect 386880 47806 386932 47812
rect 387708 47864 387760 47870
rect 387708 47806 387760 47812
rect 387984 47864 388036 47870
rect 387984 47806 388036 47812
rect 387156 4072 387208 4078
rect 387156 4014 387208 4020
rect 385960 3392 386012 3398
rect 385960 3334 386012 3340
rect 386328 3392 386380 3398
rect 386328 3334 386380 3340
rect 385972 480 386000 3334
rect 387168 480 387196 4014
rect 387720 3194 387748 47806
rect 388260 3936 388312 3942
rect 388260 3878 388312 3884
rect 387708 3188 387760 3194
rect 387708 3130 387760 3136
rect 388272 480 388300 3878
rect 389008 3466 389036 50102
rect 389088 47864 389140 47870
rect 389088 47806 389140 47812
rect 388996 3460 389048 3466
rect 388996 3402 389048 3408
rect 389100 3330 389128 47806
rect 390480 3670 390508 50102
rect 391860 3738 391888 50102
rect 392320 47870 392348 50116
rect 392308 47864 392360 47870
rect 392308 47806 392360 47812
rect 393228 47864 393280 47870
rect 393228 47806 393280 47812
rect 390652 3732 390704 3738
rect 390652 3674 390704 3680
rect 391848 3732 391900 3738
rect 391848 3674 391900 3680
rect 389456 3664 389508 3670
rect 389456 3606 389508 3612
rect 390468 3664 390520 3670
rect 390468 3606 390520 3612
rect 389088 3324 389140 3330
rect 389088 3266 389140 3272
rect 389468 480 389496 3606
rect 390664 480 390692 3674
rect 393044 3256 393096 3262
rect 393044 3198 393096 3204
rect 391848 3120 391900 3126
rect 391848 3062 391900 3068
rect 391860 480 391888 3062
rect 393056 480 393084 3198
rect 393240 3126 393268 47806
rect 393424 47530 393452 50116
rect 394542 50102 394648 50130
rect 395646 50102 396028 50130
rect 396750 50102 397408 50130
rect 393412 47524 393464 47530
rect 393412 47466 393464 47472
rect 394516 47524 394568 47530
rect 394516 47466 394568 47472
rect 394528 4078 394556 47466
rect 394516 4072 394568 4078
rect 394516 4014 394568 4020
rect 394620 3942 394648 50102
rect 394608 3936 394660 3942
rect 394608 3878 394660 3884
rect 396000 3806 396028 50102
rect 396540 4004 396592 4010
rect 396540 3946 396592 3952
rect 395344 3800 395396 3806
rect 395344 3742 395396 3748
rect 395988 3800 396040 3806
rect 395988 3742 396040 3748
rect 394240 3528 394292 3534
rect 394240 3470 394292 3476
rect 393228 3120 393280 3126
rect 393228 3062 393280 3068
rect 394252 480 394280 3470
rect 395356 480 395384 3742
rect 396552 480 396580 3946
rect 397380 3534 397408 50102
rect 397840 47598 397868 50116
rect 397828 47592 397880 47598
rect 397828 47534 397880 47540
rect 398748 47592 398800 47598
rect 398748 47534 398800 47540
rect 398760 4010 398788 47534
rect 398944 47462 398972 50116
rect 400062 50102 400168 50130
rect 401166 50102 401548 50130
rect 402178 50102 402928 50130
rect 398932 47456 398984 47462
rect 398932 47398 398984 47404
rect 400036 47456 400088 47462
rect 400036 47398 400088 47404
rect 399944 4140 399996 4146
rect 399944 4082 399996 4088
rect 398748 4004 398800 4010
rect 398748 3946 398800 3952
rect 397736 3868 397788 3874
rect 397736 3810 397788 3816
rect 397368 3528 397420 3534
rect 397368 3470 397420 3476
rect 397748 480 397776 3810
rect 398932 3596 398984 3602
rect 398932 3538 398984 3544
rect 398944 480 398972 3538
rect 399956 2122 399984 4082
rect 400048 3602 400076 47398
rect 400140 3874 400168 50102
rect 400128 3868 400180 3874
rect 400128 3810 400180 3816
rect 400036 3596 400088 3602
rect 400036 3538 400088 3544
rect 401324 3392 401376 3398
rect 401324 3334 401376 3340
rect 399956 2094 400168 2122
rect 400140 480 400168 2094
rect 401336 480 401364 3334
rect 401520 3262 401548 50102
rect 401508 3256 401560 3262
rect 401508 3198 401560 3204
rect 402520 3188 402572 3194
rect 402520 3130 402572 3136
rect 402532 480 402560 3130
rect 402900 3058 402928 50102
rect 403268 47870 403296 50116
rect 404372 47870 404400 50116
rect 405490 50102 405596 50130
rect 406594 50102 407068 50130
rect 407698 50102 408448 50130
rect 403256 47864 403308 47870
rect 403256 47806 403308 47812
rect 404268 47864 404320 47870
rect 404268 47806 404320 47812
rect 404360 47864 404412 47870
rect 404360 47806 404412 47812
rect 403624 3324 403676 3330
rect 403624 3266 403676 3272
rect 402888 3052 402940 3058
rect 402888 2994 402940 3000
rect 403636 480 403664 3266
rect 404280 2990 404308 47806
rect 405568 3466 405596 50102
rect 405648 47864 405700 47870
rect 405648 47806 405700 47812
rect 404820 3460 404872 3466
rect 404820 3402 404872 3408
rect 405556 3460 405608 3466
rect 405556 3402 405608 3408
rect 404268 2984 404320 2990
rect 404268 2926 404320 2932
rect 404832 480 404860 3402
rect 405660 3330 405688 47806
rect 407040 3670 407068 50102
rect 408420 6914 408448 50102
rect 408788 47870 408816 50116
rect 409892 47870 409920 50116
rect 411010 50102 411208 50130
rect 412114 50102 412588 50130
rect 413218 50102 413968 50130
rect 408776 47864 408828 47870
rect 408776 47806 408828 47812
rect 409788 47864 409840 47870
rect 409788 47806 409840 47812
rect 409880 47864 409932 47870
rect 409880 47806 409932 47812
rect 411076 47864 411128 47870
rect 411076 47806 411128 47812
rect 408328 6886 408448 6914
rect 407212 3732 407264 3738
rect 407212 3674 407264 3680
rect 406016 3664 406068 3670
rect 406016 3606 406068 3612
rect 407028 3664 407080 3670
rect 407028 3606 407080 3612
rect 405648 3324 405700 3330
rect 405648 3266 405700 3272
rect 406028 480 406056 3606
rect 407224 480 407252 3674
rect 408328 3194 408356 6886
rect 409604 4072 409656 4078
rect 409604 4014 409656 4020
rect 408316 3188 408368 3194
rect 408316 3130 408368 3136
rect 408408 3120 408460 3126
rect 408408 3062 408460 3068
rect 408420 480 408448 3062
rect 409616 480 409644 4014
rect 409800 3330 409828 47806
rect 411088 4146 411116 47806
rect 411076 4140 411128 4146
rect 411076 4082 411128 4088
rect 410800 3936 410852 3942
rect 410800 3878 410852 3884
rect 409788 3324 409840 3330
rect 409788 3266 409840 3272
rect 410812 480 410840 3878
rect 411180 3738 411208 50102
rect 412560 3942 412588 50102
rect 412548 3936 412600 3942
rect 412548 3878 412600 3884
rect 411904 3800 411956 3806
rect 411904 3742 411956 3748
rect 411168 3732 411220 3738
rect 411168 3674 411220 3680
rect 411916 480 411944 3742
rect 413100 3528 413152 3534
rect 413100 3470 413152 3476
rect 413112 480 413140 3470
rect 413940 3398 413968 50102
rect 414216 47462 414244 50116
rect 415228 50102 415334 50130
rect 416438 50102 416728 50130
rect 417542 50102 418108 50130
rect 414204 47456 414256 47462
rect 414204 47398 414256 47404
rect 414296 4004 414348 4010
rect 414296 3946 414348 3952
rect 413928 3392 413980 3398
rect 413928 3334 413980 3340
rect 414308 480 414336 3946
rect 415228 3534 415256 50102
rect 415308 47456 415360 47462
rect 415308 47398 415360 47404
rect 415320 3806 415348 47398
rect 416700 4078 416728 50102
rect 416688 4072 416740 4078
rect 416688 4014 416740 4020
rect 416688 3868 416740 3874
rect 416688 3810 416740 3816
rect 415308 3800 415360 3806
rect 415308 3742 415360 3748
rect 415492 3596 415544 3602
rect 415492 3538 415544 3544
rect 415216 3528 415268 3534
rect 415216 3470 415268 3476
rect 415504 480 415532 3538
rect 416700 480 416728 3810
rect 418080 3262 418108 50102
rect 418632 47870 418660 50116
rect 419736 47870 419764 50116
rect 418620 47864 418672 47870
rect 418620 47806 418672 47812
rect 419448 47864 419500 47870
rect 419448 47806 419500 47812
rect 419724 47864 419776 47870
rect 419724 47806 419776 47812
rect 420736 47864 420788 47870
rect 420736 47806 420788 47812
rect 417884 3256 417936 3262
rect 417884 3198 417936 3204
rect 418068 3256 418120 3262
rect 418068 3198 418120 3204
rect 417896 480 417924 3198
rect 419460 3058 419488 47806
rect 420748 4010 420776 47806
rect 420736 4004 420788 4010
rect 420736 3946 420788 3952
rect 420840 3602 420868 50116
rect 421958 50102 422248 50130
rect 423062 50102 423628 50130
rect 422220 3874 422248 50102
rect 422208 3868 422260 3874
rect 422208 3810 422260 3816
rect 420828 3596 420880 3602
rect 420828 3538 420880 3544
rect 422576 3460 422628 3466
rect 422576 3402 422628 3408
rect 421380 3188 421432 3194
rect 421380 3130 421432 3136
rect 418988 3052 419040 3058
rect 418988 2994 419040 3000
rect 419448 3052 419500 3058
rect 419448 2994 419500 3000
rect 419000 480 419028 2994
rect 420184 2984 420236 2990
rect 420184 2926 420236 2932
rect 420196 480 420224 2926
rect 421392 480 421420 3130
rect 422588 480 422616 3402
rect 423600 2990 423628 50102
rect 424152 47598 424180 50116
rect 424140 47592 424192 47598
rect 424140 47534 424192 47540
rect 424968 47592 425020 47598
rect 424968 47534 425020 47540
rect 424980 6914 425008 47534
rect 425256 47462 425284 50116
rect 425244 47456 425296 47462
rect 425244 47398 425296 47404
rect 424888 6886 425008 6914
rect 423772 3664 423824 3670
rect 423772 3606 423824 3612
rect 423588 2984 423640 2990
rect 423588 2926 423640 2932
rect 423784 480 423812 3606
rect 424888 3194 424916 6886
rect 426268 3466 426296 50116
rect 427386 50102 427768 50130
rect 428490 50102 429148 50130
rect 426348 47456 426400 47462
rect 426348 47398 426400 47404
rect 426256 3460 426308 3466
rect 426256 3402 426308 3408
rect 426164 3324 426216 3330
rect 426164 3266 426216 3272
rect 424876 3188 424928 3194
rect 424876 3130 424928 3136
rect 424968 3120 425020 3126
rect 424968 3062 425020 3068
rect 424980 480 425008 3062
rect 426176 480 426204 3266
rect 426360 2922 426388 47398
rect 427268 4140 427320 4146
rect 427268 4082 427320 4088
rect 426348 2916 426400 2922
rect 426348 2858 426400 2864
rect 427280 480 427308 4082
rect 427740 3670 427768 50102
rect 429120 4146 429148 50102
rect 429580 47870 429608 50116
rect 430684 47870 430712 50116
rect 429568 47864 429620 47870
rect 429568 47806 429620 47812
rect 430488 47864 430540 47870
rect 430488 47806 430540 47812
rect 430672 47864 430724 47870
rect 430672 47806 430724 47812
rect 429108 4140 429160 4146
rect 429108 4082 429160 4088
rect 430500 3942 430528 47806
rect 429660 3936 429712 3942
rect 429660 3878 429712 3884
rect 430488 3936 430540 3942
rect 430488 3878 430540 3884
rect 428464 3732 428516 3738
rect 428464 3674 428516 3680
rect 427728 3664 427780 3670
rect 427728 3606 427780 3612
rect 428476 480 428504 3674
rect 429672 480 429700 3878
rect 431788 3738 431816 50116
rect 432906 50102 433288 50130
rect 434010 50102 434668 50130
rect 431868 47864 431920 47870
rect 431868 47806 431920 47812
rect 431776 3732 431828 3738
rect 431776 3674 431828 3680
rect 430856 3392 430908 3398
rect 430856 3334 430908 3340
rect 430868 480 430896 3334
rect 431880 3330 431908 47806
rect 433260 6914 433288 50102
rect 433168 6886 433288 6914
rect 432052 3800 432104 3806
rect 432052 3742 432104 3748
rect 431868 3324 431920 3330
rect 431868 3266 431920 3272
rect 432064 480 432092 3742
rect 433168 3194 433196 6886
rect 434640 4078 434668 50102
rect 435100 47802 435128 50116
rect 436204 47870 436232 50116
rect 437230 50102 437428 50130
rect 438334 50102 438808 50130
rect 436192 47864 436244 47870
rect 436192 47806 436244 47812
rect 437296 47864 437348 47870
rect 437296 47806 437348 47812
rect 435088 47796 435140 47802
rect 435088 47738 435140 47744
rect 436008 47796 436060 47802
rect 436008 47738 436060 47744
rect 434444 4072 434496 4078
rect 434444 4014 434496 4020
rect 434628 4072 434680 4078
rect 434628 4014 434680 4020
rect 433248 3528 433300 3534
rect 433248 3470 433300 3476
rect 433156 3188 433208 3194
rect 433156 3130 433208 3136
rect 433260 480 433288 3470
rect 434456 480 434484 4014
rect 435548 3256 435600 3262
rect 435548 3198 435600 3204
rect 435560 480 435588 3198
rect 436020 2854 436048 47738
rect 437308 3806 437336 47806
rect 437296 3800 437348 3806
rect 437296 3742 437348 3748
rect 437400 3534 437428 50102
rect 437940 4004 437992 4010
rect 437940 3946 437992 3952
rect 437388 3528 437440 3534
rect 437388 3470 437440 3476
rect 436744 3052 436796 3058
rect 436744 2994 436796 3000
rect 436008 2848 436060 2854
rect 436008 2790 436060 2796
rect 436756 480 436784 2994
rect 437952 480 437980 3946
rect 438780 3058 438808 50102
rect 439424 47870 439452 50116
rect 440528 47870 440556 50116
rect 441632 47870 441660 50116
rect 442750 50102 442856 50130
rect 443854 50102 444328 50130
rect 439412 47864 439464 47870
rect 439412 47806 439464 47812
rect 440148 47864 440200 47870
rect 440148 47806 440200 47812
rect 440516 47864 440568 47870
rect 440516 47806 440568 47812
rect 441528 47864 441580 47870
rect 441528 47806 441580 47812
rect 441620 47864 441672 47870
rect 441620 47806 441672 47812
rect 439136 3596 439188 3602
rect 439136 3538 439188 3544
rect 438768 3052 438820 3058
rect 438768 2994 438820 3000
rect 439148 480 439176 3538
rect 440160 3262 440188 47806
rect 441540 4010 441568 47806
rect 441528 4004 441580 4010
rect 441528 3946 441580 3952
rect 440332 3868 440384 3874
rect 440332 3810 440384 3816
rect 440148 3256 440200 3262
rect 440148 3198 440200 3204
rect 440344 480 440372 3810
rect 442828 3602 442856 50102
rect 442908 47864 442960 47870
rect 442908 47806 442960 47812
rect 442816 3596 442868 3602
rect 442816 3538 442868 3544
rect 442632 3120 442684 3126
rect 442632 3062 442684 3068
rect 441528 2984 441580 2990
rect 441528 2926 441580 2932
rect 441540 480 441568 2926
rect 442644 480 442672 3062
rect 442920 2990 442948 47806
rect 444300 3874 444328 50102
rect 444944 47598 444972 50116
rect 446048 47870 446076 50116
rect 446036 47864 446088 47870
rect 446036 47806 446088 47812
rect 447048 47864 447100 47870
rect 447048 47806 447100 47812
rect 444932 47592 444984 47598
rect 444932 47534 444984 47540
rect 445668 47592 445720 47598
rect 445668 47534 445720 47540
rect 444288 3868 444340 3874
rect 444288 3810 444340 3816
rect 445024 3460 445076 3466
rect 445024 3402 445076 3408
rect 442908 2984 442960 2990
rect 442908 2926 442960 2932
rect 443828 2916 443880 2922
rect 443828 2858 443880 2864
rect 443840 480 443868 2858
rect 445036 480 445064 3402
rect 445680 3398 445708 47534
rect 446220 3664 446272 3670
rect 446220 3606 446272 3612
rect 445668 3392 445720 3398
rect 445668 3334 445720 3340
rect 446232 480 446260 3606
rect 447060 2990 447088 47806
rect 447152 47462 447180 50116
rect 448270 50102 448376 50130
rect 449282 50102 449848 50130
rect 447140 47456 447192 47462
rect 447140 47398 447192 47404
rect 447416 4140 447468 4146
rect 447416 4082 447468 4088
rect 447048 2984 447100 2990
rect 447048 2926 447100 2932
rect 447428 480 447456 4082
rect 448348 3670 448376 50102
rect 448428 47456 448480 47462
rect 448428 47398 448480 47404
rect 448336 3664 448388 3670
rect 448336 3606 448388 3612
rect 448440 3126 448468 47398
rect 448612 3936 448664 3942
rect 448612 3878 448664 3884
rect 448428 3120 448480 3126
rect 448428 3062 448480 3068
rect 448624 480 448652 3878
rect 449820 3482 449848 50102
rect 450372 47870 450400 50116
rect 451476 47870 451504 50116
rect 452488 50102 452594 50130
rect 453698 50102 453988 50130
rect 454802 50102 455368 50130
rect 450360 47864 450412 47870
rect 450360 47806 450412 47812
rect 451188 47864 451240 47870
rect 451188 47806 451240 47812
rect 451464 47864 451516 47870
rect 451464 47806 451516 47812
rect 451200 4146 451228 47806
rect 451188 4140 451240 4146
rect 451188 4082 451240 4088
rect 452488 3738 452516 50102
rect 452568 47864 452620 47870
rect 452568 47806 452620 47812
rect 450912 3732 450964 3738
rect 450912 3674 450964 3680
rect 452476 3732 452528 3738
rect 452476 3674 452528 3680
rect 449820 3466 449940 3482
rect 449820 3460 449952 3466
rect 449820 3454 449900 3460
rect 449900 3402 449952 3408
rect 449716 3324 449768 3330
rect 449716 3266 449768 3272
rect 449728 1714 449756 3266
rect 449728 1686 449848 1714
rect 449820 480 449848 1686
rect 450924 480 450952 3674
rect 452580 3194 452608 47806
rect 453304 4072 453356 4078
rect 453304 4014 453356 4020
rect 452108 3188 452160 3194
rect 452108 3130 452160 3136
rect 452568 3188 452620 3194
rect 452568 3130 452620 3136
rect 452120 480 452148 3130
rect 453316 480 453344 4014
rect 453960 3738 453988 50102
rect 453948 3732 454000 3738
rect 453948 3674 454000 3680
rect 455340 3194 455368 50102
rect 455892 47598 455920 50116
rect 456996 47870 457024 50116
rect 456984 47864 457036 47870
rect 456984 47806 457036 47812
rect 457996 47864 458048 47870
rect 457996 47806 458048 47812
rect 455880 47592 455932 47598
rect 455880 47534 455932 47540
rect 456708 47592 456760 47598
rect 456708 47534 456760 47540
rect 456720 4078 456748 47534
rect 456708 4072 456760 4078
rect 456708 4014 456760 4020
rect 458008 3942 458036 47806
rect 457996 3936 458048 3942
rect 457996 3878 458048 3884
rect 455696 3800 455748 3806
rect 455696 3742 455748 3748
rect 455328 3188 455380 3194
rect 455328 3130 455380 3136
rect 454500 2848 454552 2854
rect 454500 2790 454552 2796
rect 454512 480 454540 2790
rect 455708 480 455736 3742
rect 458100 3534 458128 50116
rect 459218 50102 459508 50130
rect 460322 50102 460888 50130
rect 459480 4826 459508 50102
rect 459468 4820 459520 4826
rect 459468 4762 459520 4768
rect 460388 4004 460440 4010
rect 460388 3946 460440 3952
rect 456892 3528 456944 3534
rect 456892 3470 456944 3476
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 456904 480 456932 3470
rect 459192 3256 459244 3262
rect 459192 3198 459244 3204
rect 458088 3052 458140 3058
rect 458088 2994 458140 3000
rect 458100 480 458128 2994
rect 459204 480 459232 3198
rect 460400 480 460428 3946
rect 460860 3806 460888 50102
rect 461320 47870 461348 50116
rect 461308 47864 461360 47870
rect 461308 47806 461360 47812
rect 462228 47864 462280 47870
rect 462228 47806 462280 47812
rect 460848 3800 460900 3806
rect 460848 3742 460900 3748
rect 462240 3262 462268 47806
rect 462424 47598 462452 50116
rect 463542 50102 463648 50130
rect 464646 50102 465028 50130
rect 465750 50102 466408 50130
rect 462412 47592 462464 47598
rect 462412 47534 462464 47540
rect 463620 4010 463648 50102
rect 463608 4004 463660 4010
rect 463608 3946 463660 3952
rect 463976 3868 464028 3874
rect 463976 3810 464028 3816
rect 462780 3596 462832 3602
rect 462780 3538 462832 3544
rect 462228 3256 462280 3262
rect 462228 3198 462280 3204
rect 461584 2916 461636 2922
rect 461584 2858 461636 2864
rect 461596 480 461624 2858
rect 462792 480 462820 3538
rect 463988 480 464016 3810
rect 465000 3602 465028 50102
rect 466380 5030 466408 50102
rect 466840 47870 466868 50116
rect 467944 47870 467972 50116
rect 466828 47864 466880 47870
rect 466828 47806 466880 47812
rect 467748 47864 467800 47870
rect 467748 47806 467800 47812
rect 467932 47864 467984 47870
rect 467932 47806 467984 47812
rect 466368 5024 466420 5030
rect 466368 4966 466420 4972
rect 464988 3596 465040 3602
rect 464988 3538 465040 3544
rect 465172 3392 465224 3398
rect 465172 3334 465224 3340
rect 465184 480 465212 3334
rect 467760 3126 467788 47806
rect 469048 7614 469076 50116
rect 470166 50102 470548 50130
rect 471270 50102 471928 50130
rect 469128 47864 469180 47870
rect 469128 47806 469180 47812
rect 469036 7608 469088 7614
rect 469036 7550 469088 7556
rect 468668 3664 468720 3670
rect 468668 3606 468720 3612
rect 467472 3120 467524 3126
rect 467472 3062 467524 3068
rect 467748 3120 467800 3126
rect 467748 3062 467800 3068
rect 466276 2984 466328 2990
rect 466276 2926 466328 2932
rect 466288 480 466316 2926
rect 467484 480 467512 3062
rect 468680 480 468708 3606
rect 469140 3398 469168 47806
rect 470520 3874 470548 50102
rect 471060 4140 471112 4146
rect 471060 4082 471112 4088
rect 470508 3868 470560 3874
rect 470508 3810 470560 3816
rect 469128 3392 469180 3398
rect 469128 3334 469180 3340
rect 469864 3324 469916 3330
rect 469864 3266 469916 3272
rect 469876 480 469904 3266
rect 471072 480 471100 4082
rect 471900 3330 471928 50102
rect 472268 47870 472296 50116
rect 473372 47870 473400 50116
rect 474490 50102 474688 50130
rect 475594 50102 476068 50130
rect 476698 50102 477448 50130
rect 472256 47864 472308 47870
rect 472256 47806 472308 47812
rect 473268 47864 473320 47870
rect 473268 47806 473320 47812
rect 473360 47864 473412 47870
rect 473360 47806 473412 47812
rect 474556 47864 474608 47870
rect 474556 47806 474608 47812
rect 473280 5098 473308 47806
rect 474568 11898 474596 47806
rect 474556 11892 474608 11898
rect 474556 11834 474608 11840
rect 474660 11778 474688 50102
rect 474476 11750 474688 11778
rect 473268 5092 473320 5098
rect 473268 5034 473320 5040
rect 474476 3670 474504 11750
rect 474648 11688 474700 11694
rect 474648 11630 474700 11636
rect 474660 3738 474688 11630
rect 476040 4894 476068 50102
rect 476028 4888 476080 4894
rect 476028 4830 476080 4836
rect 477420 4146 477448 50102
rect 477788 47870 477816 50116
rect 478892 47870 478920 50116
rect 480010 50102 480208 50130
rect 481114 50102 481588 50130
rect 482218 50102 482968 50130
rect 477776 47864 477828 47870
rect 477776 47806 477828 47812
rect 478788 47864 478840 47870
rect 478788 47806 478840 47812
rect 478880 47864 478932 47870
rect 478880 47806 478932 47812
rect 480076 47864 480128 47870
rect 480076 47806 480128 47812
rect 477408 4140 477460 4146
rect 477408 4082 477460 4088
rect 476948 4072 477000 4078
rect 476948 4014 477000 4020
rect 474556 3732 474608 3738
rect 474556 3674 474608 3680
rect 474648 3732 474700 3738
rect 474648 3674 474700 3680
rect 474464 3664 474516 3670
rect 474464 3606 474516 3612
rect 473452 3460 473504 3466
rect 473452 3402 473504 3408
rect 471888 3324 471940 3330
rect 471888 3266 471940 3272
rect 472256 2848 472308 2854
rect 472256 2790 472308 2796
rect 472268 480 472296 2790
rect 473464 480 473492 3402
rect 474568 480 474596 3674
rect 475752 3188 475804 3194
rect 475752 3130 475804 3136
rect 475764 480 475792 3130
rect 476960 480 476988 4014
rect 478144 3936 478196 3942
rect 478144 3878 478196 3884
rect 478156 480 478184 3878
rect 478800 3194 478828 47806
rect 480088 7682 480116 47806
rect 480076 7676 480128 7682
rect 480076 7618 480128 7624
rect 480180 3534 480208 50102
rect 480536 4820 480588 4826
rect 480536 4762 480588 4768
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 480168 3528 480220 3534
rect 480168 3470 480220 3476
rect 478788 3188 478840 3194
rect 478788 3130 478840 3136
rect 479352 480 479380 3470
rect 480548 480 480576 4762
rect 481560 4078 481588 50102
rect 482284 47592 482336 47598
rect 482284 47534 482336 47540
rect 482296 4214 482324 47534
rect 482940 4826 482968 50102
rect 483308 47870 483336 50116
rect 483296 47864 483348 47870
rect 483296 47806 483348 47812
rect 484216 47864 484268 47870
rect 484216 47806 484268 47812
rect 482928 4820 482980 4826
rect 482928 4762 482980 4768
rect 482284 4208 482336 4214
rect 482284 4150 482336 4156
rect 484032 4208 484084 4214
rect 484032 4150 484084 4156
rect 481548 4072 481600 4078
rect 481548 4014 481600 4020
rect 481732 3800 481784 3806
rect 481732 3742 481784 3748
rect 481744 480 481772 3742
rect 482836 3256 482888 3262
rect 482836 3198 482888 3204
rect 482848 480 482876 3198
rect 484044 480 484072 4150
rect 484228 3806 484256 47806
rect 484320 3942 484348 50116
rect 485438 50102 485728 50130
rect 486542 50102 487108 50130
rect 485700 4962 485728 50102
rect 485688 4956 485740 4962
rect 485688 4898 485740 4904
rect 487080 4010 487108 50102
rect 487632 47598 487660 50116
rect 488736 47598 488764 50116
rect 487620 47592 487672 47598
rect 487620 47534 487672 47540
rect 488448 47592 488500 47598
rect 488448 47534 488500 47540
rect 488724 47592 488776 47598
rect 488724 47534 488776 47540
rect 487620 5024 487672 5030
rect 487620 4966 487672 4972
rect 485228 4004 485280 4010
rect 485228 3946 485280 3952
rect 487068 4004 487120 4010
rect 487068 3946 487120 3952
rect 484308 3936 484360 3942
rect 484308 3878 484360 3884
rect 484216 3800 484268 3806
rect 484216 3742 484268 3748
rect 485240 480 485268 3946
rect 486424 3596 486476 3602
rect 486424 3538 486476 3544
rect 486436 480 486464 3538
rect 487632 480 487660 4966
rect 488460 3262 488488 47534
rect 489840 3602 489868 50116
rect 490958 50102 491248 50130
rect 491116 7608 491168 7614
rect 491116 7550 491168 7556
rect 489828 3596 489880 3602
rect 489828 3538 489880 3544
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 488448 3256 488500 3262
rect 488448 3198 488500 3204
rect 488816 3120 488868 3126
rect 488816 3062 488868 3068
rect 488828 480 488856 3062
rect 489932 480 489960 3334
rect 491128 480 491156 7550
rect 491220 3466 491248 50102
rect 492048 47326 492076 50116
rect 493152 47870 493180 50116
rect 494256 47870 494284 50116
rect 495268 50102 495374 50130
rect 496386 50102 496768 50130
rect 497490 50102 498148 50130
rect 493140 47864 493192 47870
rect 493140 47806 493192 47812
rect 493968 47864 494020 47870
rect 493968 47806 494020 47812
rect 494244 47864 494296 47870
rect 494244 47806 494296 47812
rect 492036 47320 492088 47326
rect 492036 47262 492088 47268
rect 493980 3874 494008 47806
rect 495268 47666 495296 50102
rect 495348 47864 495400 47870
rect 495348 47806 495400 47812
rect 495256 47660 495308 47666
rect 495256 47602 495308 47608
rect 494704 5092 494756 5098
rect 494704 5034 494756 5040
rect 492312 3868 492364 3874
rect 492312 3810 492364 3816
rect 493968 3868 494020 3874
rect 493968 3810 494020 3816
rect 491208 3460 491260 3466
rect 491208 3402 491260 3408
rect 492324 480 492352 3810
rect 493508 3324 493560 3330
rect 493508 3266 493560 3272
rect 493520 480 493548 3266
rect 494716 480 494744 5034
rect 495360 3058 495388 47806
rect 496740 3738 496768 50102
rect 497464 47320 497516 47326
rect 497464 47262 497516 47268
rect 497476 7614 497504 47262
rect 497464 7608 497516 7614
rect 497464 7550 497516 7556
rect 495900 3732 495952 3738
rect 495900 3674 495952 3680
rect 496728 3732 496780 3738
rect 496728 3674 496780 3680
rect 495348 3052 495400 3058
rect 495348 2994 495400 3000
rect 495912 480 495940 3674
rect 498120 3670 498148 50102
rect 498580 47734 498608 50116
rect 499684 47870 499712 50116
rect 500802 50102 500908 50130
rect 501906 50102 502288 50130
rect 503010 50102 503668 50130
rect 499672 47864 499724 47870
rect 499672 47806 499724 47812
rect 500776 47864 500828 47870
rect 500776 47806 500828 47812
rect 498568 47728 498620 47734
rect 498568 47670 498620 47676
rect 498200 4888 498252 4894
rect 498200 4830 498252 4836
rect 497096 3664 497148 3670
rect 497096 3606 497148 3612
rect 498108 3664 498160 3670
rect 498108 3606 498160 3612
rect 497108 480 497136 3606
rect 498212 480 498240 4830
rect 499396 4140 499448 4146
rect 499396 4082 499448 4088
rect 499408 480 499436 4082
rect 500592 3188 500644 3194
rect 500592 3130 500644 3136
rect 500604 480 500632 3130
rect 500788 3126 500816 47806
rect 500880 3398 500908 50102
rect 501788 7676 501840 7682
rect 501788 7618 501840 7624
rect 500868 3392 500920 3398
rect 500868 3334 500920 3340
rect 500776 3120 500828 3126
rect 500776 3062 500828 3068
rect 501800 480 501828 7618
rect 502260 5098 502288 50102
rect 502984 47728 503036 47734
rect 502984 47670 503036 47676
rect 502996 5234 503024 47670
rect 502984 5228 503036 5234
rect 502984 5170 503036 5176
rect 502248 5092 502300 5098
rect 502248 5034 502300 5040
rect 502984 3528 503036 3534
rect 502984 3470 503036 3476
rect 502996 480 503024 3470
rect 503640 3330 503668 50102
rect 504100 47870 504128 50116
rect 504088 47864 504140 47870
rect 504088 47806 504140 47812
rect 505008 47864 505060 47870
rect 505008 47806 505060 47812
rect 504364 47660 504416 47666
rect 504364 47602 504416 47608
rect 504376 7682 504404 47602
rect 504364 7676 504416 7682
rect 504364 7618 504416 7624
rect 505020 4146 505048 47806
rect 505204 47666 505232 50116
rect 506322 50102 506428 50130
rect 507426 50102 507808 50130
rect 505192 47660 505244 47666
rect 505192 47602 505244 47608
rect 505376 4820 505428 4826
rect 505376 4762 505428 4768
rect 505008 4140 505060 4146
rect 505008 4082 505060 4088
rect 504180 4072 504232 4078
rect 504180 4014 504232 4020
rect 503628 3324 503680 3330
rect 503628 3266 503680 3272
rect 504192 480 504220 4014
rect 505388 480 505416 4762
rect 506400 3534 506428 50102
rect 507780 3942 507808 50102
rect 508424 47870 508452 50116
rect 508412 47864 508464 47870
rect 508412 47806 508464 47812
rect 509148 47864 509200 47870
rect 509148 47806 509200 47812
rect 509160 5166 509188 47806
rect 509528 47734 509556 50116
rect 510632 47870 510660 50116
rect 511750 50102 511856 50130
rect 512854 50102 513328 50130
rect 510620 47864 510672 47870
rect 510620 47806 510672 47812
rect 509516 47728 509568 47734
rect 509516 47670 509568 47676
rect 510528 47728 510580 47734
rect 510528 47670 510580 47676
rect 509148 5160 509200 5166
rect 509148 5102 509200 5108
rect 508872 4956 508924 4962
rect 508872 4898 508924 4904
rect 507676 3936 507728 3942
rect 507676 3878 507728 3884
rect 507768 3936 507820 3942
rect 507768 3878 507820 3884
rect 506480 3800 506532 3806
rect 506480 3742 506532 3748
rect 506388 3528 506440 3534
rect 506388 3470 506440 3476
rect 506492 480 506520 3742
rect 507688 480 507716 3878
rect 508884 480 508912 4898
rect 510540 4078 510568 47670
rect 511828 4894 511856 50102
rect 511908 47864 511960 47870
rect 511908 47806 511960 47812
rect 511816 4888 511868 4894
rect 511816 4830 511868 4836
rect 510528 4072 510580 4078
rect 510528 4014 510580 4020
rect 510068 4004 510120 4010
rect 510068 3946 510120 3952
rect 510080 480 510108 3946
rect 511920 3262 511948 47806
rect 512092 47592 512144 47598
rect 512092 47534 512144 47540
rect 511264 3256 511316 3262
rect 511264 3198 511316 3204
rect 511908 3256 511960 3262
rect 511908 3198 511960 3204
rect 511276 480 511304 3198
rect 512104 490 512132 47534
rect 513300 3806 513328 50102
rect 513944 47870 513972 50116
rect 515048 47870 515076 50116
rect 516152 47870 516180 50116
rect 517270 50102 517376 50130
rect 518374 50102 518848 50130
rect 513932 47864 513984 47870
rect 513932 47806 513984 47812
rect 514668 47864 514720 47870
rect 514668 47806 514720 47812
rect 515036 47864 515088 47870
rect 515036 47806 515088 47812
rect 516048 47864 516100 47870
rect 516048 47806 516100 47812
rect 516140 47864 516192 47870
rect 516140 47806 516192 47812
rect 514680 4010 514708 47806
rect 515404 47660 515456 47666
rect 515404 47602 515456 47608
rect 515416 7750 515444 47602
rect 515404 7744 515456 7750
rect 515404 7686 515456 7692
rect 516060 7614 516088 47806
rect 515956 7608 516008 7614
rect 515956 7550 516008 7556
rect 516048 7608 516100 7614
rect 516048 7550 516100 7556
rect 514668 4004 514720 4010
rect 514668 3946 514720 3952
rect 513288 3800 513340 3806
rect 513288 3742 513340 3748
rect 513564 3596 513616 3602
rect 513564 3538 513616 3544
rect 512288 598 512500 626
rect 512288 490 512316 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512104 462 512316 490
rect 512472 480 512500 598
rect 513576 480 513604 3538
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 514772 480 514800 3402
rect 515968 480 515996 7550
rect 517152 3868 517204 3874
rect 517152 3810 517204 3816
rect 517164 480 517192 3810
rect 517348 3466 517376 50102
rect 517428 47864 517480 47870
rect 517428 47806 517480 47812
rect 517336 3460 517388 3466
rect 517336 3402 517388 3408
rect 517440 3194 517468 47806
rect 518820 5030 518848 50102
rect 519372 47870 519400 50116
rect 520476 47870 520504 50116
rect 521488 50102 521594 50130
rect 522698 50102 522988 50130
rect 523802 50102 524368 50130
rect 519360 47864 519412 47870
rect 519360 47806 519412 47812
rect 520188 47864 520240 47870
rect 520188 47806 520240 47812
rect 520464 47864 520516 47870
rect 520464 47806 520516 47812
rect 519544 7676 519596 7682
rect 519544 7618 519596 7624
rect 518808 5024 518860 5030
rect 518808 4966 518860 4972
rect 517428 3188 517480 3194
rect 517428 3130 517480 3136
rect 518348 3052 518400 3058
rect 518348 2994 518400 3000
rect 518360 480 518388 2994
rect 519556 480 519584 7618
rect 520200 3602 520228 47806
rect 521488 4826 521516 50102
rect 521568 47864 521620 47870
rect 521568 47806 521620 47812
rect 521476 4820 521528 4826
rect 521476 4762 521528 4768
rect 521580 3874 521608 47806
rect 521568 3868 521620 3874
rect 521568 3810 521620 3816
rect 520740 3732 520792 3738
rect 520740 3674 520792 3680
rect 520188 3596 520240 3602
rect 520188 3538 520240 3544
rect 520752 480 520780 3674
rect 522960 3670 522988 50102
rect 523040 5228 523092 5234
rect 523040 5170 523092 5176
rect 521844 3664 521896 3670
rect 521844 3606 521896 3612
rect 522948 3664 523000 3670
rect 522948 3606 523000 3612
rect 521856 480 521884 3606
rect 523052 480 523080 5170
rect 524236 3120 524288 3126
rect 524236 3062 524288 3068
rect 524248 480 524276 3062
rect 524340 2854 524368 50102
rect 524892 47870 524920 50116
rect 525996 47870 526024 50116
rect 524880 47864 524932 47870
rect 524880 47806 524932 47812
rect 525708 47864 525760 47870
rect 525708 47806 525760 47812
rect 525984 47864 526036 47870
rect 525984 47806 526036 47812
rect 526996 47864 527048 47870
rect 526996 47806 527048 47812
rect 525720 4962 525748 47806
rect 526628 5092 526680 5098
rect 526628 5034 526680 5040
rect 525708 4956 525760 4962
rect 525708 4898 525760 4904
rect 525432 3392 525484 3398
rect 525432 3334 525484 3340
rect 524328 2848 524380 2854
rect 524328 2790 524380 2796
rect 525444 480 525472 3334
rect 526640 480 526668 5034
rect 527008 3738 527036 47806
rect 526996 3732 527048 3738
rect 526996 3674 527048 3680
rect 527100 3398 527128 50116
rect 528204 47734 528232 50116
rect 529322 50102 529888 50130
rect 528192 47728 528244 47734
rect 528192 47670 528244 47676
rect 529860 4146 529888 50102
rect 530412 47870 530440 50116
rect 531424 48006 531452 50116
rect 532542 50102 532648 50130
rect 533646 50102 534028 50130
rect 531412 48000 531464 48006
rect 531412 47942 531464 47948
rect 530400 47864 530452 47870
rect 530400 47806 530452 47812
rect 531228 47864 531280 47870
rect 531228 47806 531280 47812
rect 530124 7744 530176 7750
rect 530124 7686 530176 7692
rect 529020 4140 529072 4146
rect 529020 4082 529072 4088
rect 529848 4140 529900 4146
rect 529848 4082 529900 4088
rect 527088 3392 527140 3398
rect 527088 3334 527140 3340
rect 527824 3324 527876 3330
rect 527824 3266 527876 3272
rect 527836 480 527864 3266
rect 529032 480 529060 4082
rect 530136 480 530164 7686
rect 531240 2922 531268 47806
rect 532516 3936 532568 3942
rect 532516 3878 532568 3884
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531228 2916 531280 2922
rect 531228 2858 531280 2864
rect 531332 480 531360 3470
rect 532528 480 532556 3878
rect 532620 3330 532648 50102
rect 533712 5160 533764 5166
rect 533712 5102 533764 5108
rect 532608 3324 532660 3330
rect 532608 3266 532660 3272
rect 533724 480 533752 5102
rect 534000 2990 534028 50102
rect 534736 47802 534764 50116
rect 535840 47870 535868 50116
rect 536944 48006 536972 50116
rect 536932 48000 536984 48006
rect 536932 47942 536984 47948
rect 535828 47864 535880 47870
rect 535828 47806 535880 47812
rect 536748 47864 536800 47870
rect 536748 47806 536800 47812
rect 534724 47796 534776 47802
rect 534724 47738 534776 47744
rect 534908 4072 534960 4078
rect 534908 4014 534960 4020
rect 533988 2984 534040 2990
rect 533988 2926 534040 2932
rect 534920 480 534948 4014
rect 536760 3262 536788 47806
rect 538048 47802 538076 50116
rect 539166 50102 539548 50130
rect 540270 50102 540928 50130
rect 538128 48000 538180 48006
rect 538128 47942 538180 47948
rect 538036 47796 538088 47802
rect 538036 47738 538088 47744
rect 537208 4888 537260 4894
rect 537208 4830 537260 4836
rect 536104 3256 536156 3262
rect 536104 3198 536156 3204
rect 536748 3256 536800 3262
rect 536748 3198 536800 3204
rect 536116 480 536144 3198
rect 537220 480 537248 4830
rect 538140 3058 538168 47942
rect 539520 3942 539548 50102
rect 540796 7608 540848 7614
rect 540796 7550 540848 7556
rect 539600 4004 539652 4010
rect 539600 3946 539652 3952
rect 539508 3936 539560 3942
rect 539508 3878 539560 3884
rect 538404 3800 538456 3806
rect 538404 3742 538456 3748
rect 538128 3052 538180 3058
rect 538128 2994 538180 3000
rect 538416 480 538444 3742
rect 539612 480 539640 3946
rect 540808 480 540836 7550
rect 540900 3126 540928 50102
rect 541360 47666 541388 50116
rect 541348 47660 541400 47666
rect 541348 47602 541400 47608
rect 542464 47326 542492 50116
rect 543490 50102 543596 50130
rect 544594 50102 545068 50130
rect 545698 50102 546448 50130
rect 542452 47320 542504 47326
rect 542452 47262 542504 47268
rect 543568 3534 543596 50102
rect 543648 47320 543700 47326
rect 543648 47262 543700 47268
rect 543660 4078 543688 47262
rect 544384 5024 544436 5030
rect 544384 4966 544436 4972
rect 543648 4072 543700 4078
rect 543648 4014 543700 4020
rect 543556 3528 543608 3534
rect 543556 3470 543608 3476
rect 543188 3460 543240 3466
rect 543188 3402 543240 3408
rect 541992 3188 542044 3194
rect 541992 3130 542044 3136
rect 540888 3120 540940 3126
rect 540888 3062 540940 3068
rect 542004 480 542032 3130
rect 543200 480 543228 3402
rect 544396 480 544424 4966
rect 545040 3806 545068 50102
rect 546420 4010 546448 50102
rect 546788 48006 546816 50116
rect 547892 48006 547920 50116
rect 549010 50102 549208 50130
rect 550114 50102 550588 50130
rect 551218 50102 551968 50130
rect 546776 48000 546828 48006
rect 546776 47942 546828 47948
rect 547788 48000 547840 48006
rect 547788 47942 547840 47948
rect 547880 48000 547932 48006
rect 547880 47942 547932 47948
rect 549076 48000 549128 48006
rect 549076 47942 549128 47948
rect 546408 4004 546460 4010
rect 546408 3946 546460 3952
rect 546684 3868 546736 3874
rect 546684 3810 546736 3816
rect 545028 3800 545080 3806
rect 545028 3742 545080 3748
rect 545488 3596 545540 3602
rect 545488 3538 545540 3544
rect 545500 480 545528 3538
rect 546696 480 546724 3810
rect 547800 3194 547828 47942
rect 547880 4820 547932 4826
rect 547880 4762 547932 4768
rect 547788 3188 547840 3194
rect 547788 3130 547840 3136
rect 547892 480 547920 4762
rect 549088 3874 549116 47942
rect 549076 3868 549128 3874
rect 549076 3810 549128 3816
rect 549076 3664 549128 3670
rect 549076 3606 549128 3612
rect 549088 480 549116 3606
rect 549180 3602 549208 50102
rect 550560 3670 550588 50102
rect 551468 4956 551520 4962
rect 551468 4898 551520 4904
rect 550548 3664 550600 3670
rect 550548 3606 550600 3612
rect 549168 3596 549220 3602
rect 549168 3538 549220 3544
rect 550272 2848 550324 2854
rect 550272 2790 550324 2796
rect 550284 480 550312 2790
rect 551480 480 551508 4898
rect 551940 3466 551968 50102
rect 552308 47734 552336 50116
rect 552296 47728 552348 47734
rect 552296 47670 552348 47676
rect 553308 47728 553360 47734
rect 553308 47670 553360 47676
rect 553320 3738 553348 47670
rect 553412 47598 553440 50116
rect 553400 47592 553452 47598
rect 553400 47534 553452 47540
rect 554780 47524 554832 47530
rect 554780 47466 554832 47472
rect 554792 16574 554820 47466
rect 554792 16546 555004 16574
rect 552664 3732 552716 3738
rect 552664 3674 552716 3680
rect 553308 3732 553360 3738
rect 553308 3674 553360 3680
rect 551928 3460 551980 3466
rect 551928 3402 551980 3408
rect 552676 480 552704 3674
rect 553768 3392 553820 3398
rect 553768 3334 553820 3340
rect 553780 480 553808 3334
rect 554976 480 555004 16546
rect 556816 6866 556844 669287
rect 556896 668840 556948 668846
rect 556896 668782 556948 668788
rect 556908 471986 556936 668782
rect 557000 592006 557028 671706
rect 558182 669488 558238 669497
rect 558182 669423 558238 669432
rect 556988 592000 557040 592006
rect 556988 591942 557040 591948
rect 556896 471980 556948 471986
rect 556896 471922 556948 471928
rect 557540 47932 557592 47938
rect 557540 47874 557592 47880
rect 557552 16574 557580 47874
rect 558196 33114 558224 669423
rect 558288 179382 558316 672386
rect 565268 671900 565320 671906
rect 565268 671842 565320 671848
rect 561036 671424 561088 671430
rect 561036 671366 561088 671372
rect 558368 669928 558420 669934
rect 558368 669870 558420 669876
rect 558380 458182 558408 669870
rect 560944 669452 560996 669458
rect 560944 669394 560996 669400
rect 558368 458176 558420 458182
rect 558368 458118 558420 458124
rect 558276 179376 558328 179382
rect 558276 179318 558328 179324
rect 560956 60722 560984 669394
rect 561048 405686 561076 671366
rect 565176 671220 565228 671226
rect 565176 671162 565228 671168
rect 562508 670200 562560 670206
rect 562508 670142 562560 670148
rect 561128 669996 561180 670002
rect 561128 669938 561180 669944
rect 561140 511970 561168 669938
rect 562416 669724 562468 669730
rect 562416 669666 562468 669672
rect 562324 667956 562376 667962
rect 562324 667898 562376 667904
rect 561128 511964 561180 511970
rect 561128 511906 561180 511912
rect 561036 405680 561088 405686
rect 561036 405622 561088 405628
rect 560944 60716 560996 60722
rect 560944 60658 560996 60664
rect 560944 47864 560996 47870
rect 560944 47806 560996 47812
rect 558184 33108 558236 33114
rect 558184 33050 558236 33056
rect 557552 16546 558592 16574
rect 556804 6860 556856 6866
rect 556804 6802 556856 6808
rect 556160 4140 556212 4146
rect 556160 4082 556212 4088
rect 556172 480 556200 4082
rect 557356 2916 557408 2922
rect 557356 2858 557408 2864
rect 557368 480 557396 2858
rect 558564 480 558592 16546
rect 560956 5574 560984 47806
rect 562336 20670 562364 667898
rect 562428 353258 562456 669666
rect 562520 564398 562548 670142
rect 565084 668092 565136 668098
rect 565084 668034 565136 668040
rect 562508 564392 562560 564398
rect 562508 564334 562560 564340
rect 562416 353252 562468 353258
rect 562416 353194 562468 353200
rect 565096 113150 565124 668034
rect 565188 299470 565216 671162
rect 565280 618254 565308 671842
rect 566556 669656 566608 669662
rect 566462 669624 566518 669633
rect 566556 669598 566608 669604
rect 566462 669559 566518 669568
rect 565268 618248 565320 618254
rect 565268 618190 565320 618196
rect 565176 299464 565228 299470
rect 565176 299406 565228 299412
rect 565084 113144 565136 113150
rect 565084 113086 565136 113092
rect 564532 47796 564584 47802
rect 564532 47738 564584 47744
rect 562324 20664 562376 20670
rect 562324 20606 562376 20612
rect 564544 16574 564572 47738
rect 566476 46918 566504 669559
rect 566568 259418 566596 669598
rect 566660 431934 566688 672998
rect 576308 672988 576360 672994
rect 576308 672930 576360 672936
rect 571984 672852 572036 672858
rect 571984 672794 572036 672800
rect 570604 672580 570656 672586
rect 570604 672522 570656 672528
rect 569316 672240 569368 672246
rect 569316 672182 569368 672188
rect 569224 670744 569276 670750
rect 569224 670686 569276 670692
rect 566740 670540 566792 670546
rect 566740 670482 566792 670488
rect 566752 644434 566780 670482
rect 566740 644428 566792 644434
rect 566740 644370 566792 644376
rect 566648 431928 566700 431934
rect 566648 431870 566700 431876
rect 566556 259412 566608 259418
rect 566556 259354 566608 259360
rect 569236 86970 569264 670686
rect 569328 193186 569356 672182
rect 570616 273222 570644 672522
rect 571996 313274 572024 672794
rect 572076 672784 572128 672790
rect 572076 672726 572128 672732
rect 572088 325650 572116 672726
rect 573456 672376 573508 672382
rect 573456 672318 573508 672324
rect 573364 670812 573416 670818
rect 573364 670754 573416 670760
rect 572076 325644 572128 325650
rect 572076 325586 572128 325592
rect 571984 313268 572036 313274
rect 571984 313210 572036 313216
rect 570604 273216 570656 273222
rect 570604 273158 570656 273164
rect 569316 193180 569368 193186
rect 569316 193122 569368 193128
rect 573376 126954 573404 670754
rect 573468 233238 573496 672318
rect 576122 670712 576178 670721
rect 576122 670647 576178 670656
rect 574928 670472 574980 670478
rect 574928 670414 574980 670420
rect 574836 669520 574888 669526
rect 574836 669462 574888 669468
rect 574744 668160 574796 668166
rect 574744 668102 574796 668108
rect 573456 233232 573508 233238
rect 573456 233174 573508 233180
rect 574756 153202 574784 668102
rect 574848 167006 574876 669462
rect 574940 632058 574968 670414
rect 574928 632052 574980 632058
rect 574928 631994 574980 632000
rect 574836 167000 574888 167006
rect 574836 166942 574888 166948
rect 574744 153196 574796 153202
rect 574744 153138 574796 153144
rect 573364 126948 573416 126954
rect 573364 126890 573416 126896
rect 569224 86964 569276 86970
rect 569224 86906 569276 86912
rect 576136 73166 576164 670647
rect 576216 669588 576268 669594
rect 576216 669530 576268 669536
rect 576228 245614 576256 669530
rect 576320 365702 576348 672930
rect 578884 672308 578936 672314
rect 578884 672250 578936 672256
rect 576308 365696 576360 365702
rect 576308 365638 576360 365644
rect 576216 245608 576268 245614
rect 576216 245550 576268 245556
rect 578896 219065 578924 672250
rect 580172 671832 580224 671838
rect 580172 671774 580224 671780
rect 580184 670721 580212 671774
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580356 670676 580408 670682
rect 580356 670618 580408 670624
rect 580264 669384 580316 669390
rect 580264 669326 580316 669332
rect 578976 668500 579028 668506
rect 578976 668442 579028 668448
rect 578988 378457 579016 668442
rect 580172 644428 580224 644434
rect 580172 644370 580224 644376
rect 580184 644065 580212 644370
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 579712 632052 579764 632058
rect 579712 631994 579764 632000
rect 579724 630873 579752 631994
rect 579710 630864 579766 630873
rect 579710 630799 579766 630808
rect 579804 618248 579856 618254
rect 579804 618190 579856 618196
rect 579816 617545 579844 618190
rect 579802 617536 579858 617545
rect 579802 617471 579858 617480
rect 580172 592000 580224 592006
rect 580172 591942 580224 591948
rect 580184 591025 580212 591942
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580172 578196 580224 578202
rect 580172 578138 580224 578144
rect 580184 577697 580212 578138
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580172 525768 580224 525774
rect 580172 525710 580224 525716
rect 580184 524521 580212 525710
rect 580170 524512 580226 524521
rect 580170 524447 580226 524456
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 578974 378448 579030 378457
rect 578974 378383 579030 378392
rect 579988 365696 580040 365702
rect 579988 365638 580040 365644
rect 580000 365129 580028 365638
rect 579986 365120 580042 365129
rect 579986 365055 580042 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 579620 259412 579672 259418
rect 579620 259354 579672 259360
rect 579632 258913 579660 259354
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 578882 219056 578938 219065
rect 578882 218991 578938 219000
rect 579896 206984 579948 206990
rect 579896 206926 579948 206932
rect 579908 205737 579936 206926
rect 579894 205728 579950 205737
rect 579894 205663 579950 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579620 153196 579672 153202
rect 579620 153138 579672 153144
rect 579632 152697 579660 153138
rect 579618 152688 579674 152697
rect 579618 152623 579674 152632
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580276 99521 580304 669326
rect 580368 139369 580396 670618
rect 580448 669792 580500 669798
rect 580448 669734 580500 669740
rect 580460 418305 580488 669734
rect 580446 418296 580502 418305
rect 580446 418231 580502 418240
rect 580354 139360 580410 139369
rect 580354 139295 580410 139304
rect 580262 99512 580318 99521
rect 580262 99447 580318 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 576124 73160 576176 73166
rect 576124 73102 576176 73108
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 568580 47660 568632 47666
rect 568580 47602 568632 47608
rect 566464 46912 566516 46918
rect 566464 46854 566516 46860
rect 568592 16574 568620 47602
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 564544 16546 565216 16574
rect 568592 16546 568712 16574
rect 560944 5568 560996 5574
rect 560944 5510 560996 5516
rect 562048 5568 562100 5574
rect 562048 5510 562100 5516
rect 559748 3324 559800 3330
rect 559748 3266 559800 3272
rect 559760 480 559788 3266
rect 560852 2984 560904 2990
rect 560852 2926 560904 2932
rect 560864 480 560892 2926
rect 562060 480 562088 5510
rect 563244 3256 563296 3262
rect 563244 3198 563296 3204
rect 563256 480 563284 3198
rect 564440 3052 564492 3058
rect 564440 2994 564492 3000
rect 564452 480 564480 2994
rect 565188 490 565216 16546
rect 566832 3936 566884 3942
rect 566832 3878 566884 3884
rect 565464 598 565676 626
rect 565464 490 565492 598
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 462 565492 490
rect 565648 480 565676 598
rect 566844 480 566872 3878
rect 568028 3120 568080 3126
rect 568028 3062 568080 3068
rect 568040 480 568068 3062
rect 568684 490 568712 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 570328 4072 570380 4078
rect 570328 4014 570380 4020
rect 568960 598 569172 626
rect 568960 490 568988 598
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 462 568988 490
rect 569144 480 569172 598
rect 570340 480 570368 4014
rect 573916 4004 573968 4010
rect 573916 3946 573968 3952
rect 572720 3800 572772 3806
rect 572720 3742 572772 3748
rect 571524 3528 571576 3534
rect 571524 3470 571576 3476
rect 571536 480 571564 3470
rect 572732 480 572760 3742
rect 573928 480 573956 3946
rect 576308 3868 576360 3874
rect 576308 3810 576360 3816
rect 575112 3188 575164 3194
rect 575112 3130 575164 3136
rect 575124 480 575152 3130
rect 576320 480 576348 3810
rect 582196 3732 582248 3738
rect 582196 3674 582248 3680
rect 578608 3664 578660 3670
rect 578608 3606 578660 3612
rect 577412 3596 577464 3602
rect 577412 3538 577464 3544
rect 577424 480 577452 3538
rect 578620 480 578648 3606
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3674
rect 583392 3052 583444 3058
rect 583392 2994 583444 3000
rect 583404 480 583432 2994
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3054 671200 3110 671256
rect 3238 658180 3240 658200
rect 3240 658180 3292 658200
rect 3292 658180 3294 658200
rect 3238 658144 3294 658180
rect 3330 632032 3386 632088
rect 2962 619112 3018 619168
rect 2870 606056 2926 606112
rect 3146 579944 3202 580000
rect 3330 553832 3386 553888
rect 3238 527856 3294 527912
rect 2778 514800 2834 514856
rect 3330 501744 3386 501800
rect 3330 475632 3386 475688
rect 2778 462576 2834 462632
rect 2962 449556 2964 449576
rect 2964 449556 3016 449576
rect 3016 449556 3018 449576
rect 2962 449520 3018 449556
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 3330 371320 3386 371376
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 2962 345344 3018 345400
rect 3238 319232 3294 319288
rect 3330 306212 3332 306232
rect 3332 306212 3384 306232
rect 3384 306212 3386 306232
rect 3330 306176 3386 306212
rect 3238 267144 3294 267200
rect 3330 254088 3386 254144
rect 2778 241068 2780 241088
rect 2780 241068 2832 241088
rect 2832 241068 2834 241088
rect 2778 241032 2834 241068
rect 3330 214920 3386 214976
rect 3330 201864 3386 201920
rect 3330 162832 3386 162888
rect 2778 136720 2834 136776
rect 2962 110608 3018 110664
rect 3238 97552 3294 97608
rect 3054 58520 3110 58576
rect 2778 32408 2834 32464
rect 3882 566888 3938 566944
rect 3790 397432 3846 397488
rect 3698 293120 3754 293176
rect 3606 188808 3662 188864
rect 3606 149776 3662 149832
rect 6182 670792 6238 670848
rect 3514 84632 3570 84688
rect 3514 71612 3516 71632
rect 3516 71612 3568 71632
rect 3568 71612 3570 71632
rect 3514 71576 3570 71612
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 11702 672424 11758 672480
rect 10322 672152 10378 672208
rect 8942 670928 8998 670984
rect 13082 672288 13138 672344
rect 35070 670656 35126 670712
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 518714 672424 518770 672480
rect 532790 672288 532846 672344
rect 523406 670928 523462 670984
rect 546866 672152 546922 672208
rect 537482 670792 537538 670848
rect 30654 669568 30710 669624
rect 16486 669432 16542 669488
rect 21270 669432 21326 669488
rect 556802 669296 556858 669352
rect 558182 669432 558238 669488
rect 566462 669568 566518 669624
rect 576122 670656 576178 670712
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 579710 630808 579766 630864
rect 579802 617480 579858 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 537784 580226 537840
rect 580170 524456 580226 524512
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 431568 580226 431624
rect 580170 404912 580226 404968
rect 578974 378392 579030 378448
rect 579986 365064 580042 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 579618 258848 579674 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 578882 219000 578938 219056
rect 579894 205672 579950 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 579618 152632 579674 152688
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580446 418240 580502 418296
rect 580354 139304 580410 139360
rect 580262 99456 580318 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 11697 672482 11763 672485
rect 518709 672482 518775 672485
rect 11697 672480 518775 672482
rect 11697 672424 11702 672480
rect 11758 672424 518714 672480
rect 518770 672424 518775 672480
rect 11697 672422 518775 672424
rect 11697 672419 11763 672422
rect 518709 672419 518775 672422
rect 13077 672346 13143 672349
rect 532785 672346 532851 672349
rect 13077 672344 532851 672346
rect 13077 672288 13082 672344
rect 13138 672288 532790 672344
rect 532846 672288 532851 672344
rect 13077 672286 532851 672288
rect 13077 672283 13143 672286
rect 532785 672283 532851 672286
rect 10317 672210 10383 672213
rect 546861 672210 546927 672213
rect 10317 672208 546927 672210
rect 10317 672152 10322 672208
rect 10378 672152 546866 672208
rect 546922 672152 546927 672208
rect 10317 672150 546927 672152
rect 10317 672147 10383 672150
rect 546861 672147 546927 672150
rect -960 671258 480 671348
rect 3049 671258 3115 671261
rect -960 671256 3115 671258
rect -960 671200 3054 671256
rect 3110 671200 3115 671256
rect -960 671198 3115 671200
rect -960 671108 480 671198
rect 3049 671195 3115 671198
rect 8937 670986 9003 670989
rect 523401 670986 523467 670989
rect 8937 670984 523467 670986
rect 8937 670928 8942 670984
rect 8998 670928 523406 670984
rect 523462 670928 523467 670984
rect 8937 670926 523467 670928
rect 8937 670923 9003 670926
rect 523401 670923 523467 670926
rect 6177 670850 6243 670853
rect 537477 670850 537543 670853
rect 6177 670848 537543 670850
rect 6177 670792 6182 670848
rect 6238 670792 537482 670848
rect 537538 670792 537543 670848
rect 6177 670790 537543 670792
rect 6177 670787 6243 670790
rect 537477 670787 537543 670790
rect 35065 670714 35131 670717
rect 576117 670714 576183 670717
rect 35065 670712 576183 670714
rect 35065 670656 35070 670712
rect 35126 670656 576122 670712
rect 576178 670656 576183 670712
rect 35065 670654 576183 670656
rect 35065 670651 35131 670654
rect 576117 670651 576183 670654
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 30649 669626 30715 669629
rect 566457 669626 566523 669629
rect 30649 669624 566523 669626
rect 30649 669568 30654 669624
rect 30710 669568 566462 669624
rect 566518 669568 566523 669624
rect 30649 669566 566523 669568
rect 30649 669563 30715 669566
rect 566457 669563 566523 669566
rect 16481 669490 16547 669493
rect 21265 669490 21331 669493
rect 558177 669490 558243 669493
rect 16481 669488 16590 669490
rect 16481 669432 16486 669488
rect 16542 669432 16590 669488
rect 16481 669427 16590 669432
rect 21265 669488 558243 669490
rect 21265 669432 21270 669488
rect 21326 669432 558182 669488
rect 558238 669432 558243 669488
rect 21265 669430 558243 669432
rect 21265 669427 21331 669430
rect 558177 669427 558243 669430
rect 16530 669354 16590 669427
rect 556797 669354 556863 669357
rect 16530 669352 556863 669354
rect 16530 669296 556802 669352
rect 556858 669296 556863 669352
rect 16530 669294 556863 669296
rect 556797 669291 556863 669294
rect -960 658202 480 658292
rect 3233 658202 3299 658205
rect -960 658200 3299 658202
rect -960 658144 3238 658200
rect 3294 658144 3299 658200
rect -960 658142 3299 658144
rect -960 658052 480 658142
rect 3233 658139 3299 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3325 632090 3391 632093
rect -960 632088 3391 632090
rect -960 632032 3330 632088
rect 3386 632032 3391 632088
rect -960 632030 3391 632032
rect -960 631940 480 632030
rect 3325 632027 3391 632030
rect 579705 630866 579771 630869
rect 583520 630866 584960 630956
rect 579705 630864 584960 630866
rect 579705 630808 579710 630864
rect 579766 630808 584960 630864
rect 579705 630806 584960 630808
rect 579705 630803 579771 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2957 619170 3023 619173
rect -960 619168 3023 619170
rect -960 619112 2962 619168
rect 3018 619112 3023 619168
rect -960 619110 3023 619112
rect -960 619020 480 619110
rect 2957 619107 3023 619110
rect 579797 617538 579863 617541
rect 583520 617538 584960 617628
rect 579797 617536 584960 617538
rect 579797 617480 579802 617536
rect 579858 617480 584960 617536
rect 579797 617478 584960 617480
rect 579797 617475 579863 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 2865 606114 2931 606117
rect -960 606112 2931 606114
rect -960 606056 2870 606112
rect 2926 606056 2931 606112
rect -960 606054 2931 606056
rect -960 605964 480 606054
rect 2865 606051 2931 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3877 566946 3943 566949
rect -960 566944 3943 566946
rect -960 566888 3882 566944
rect 3938 566888 3943 566944
rect -960 566886 3943 566888
rect -960 566796 480 566886
rect 3877 566883 3943 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3233 527914 3299 527917
rect -960 527912 3299 527914
rect -960 527856 3238 527912
rect 3294 527856 3299 527912
rect -960 527854 3299 527856
rect -960 527764 480 527854
rect 3233 527851 3299 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 2957 449578 3023 449581
rect -960 449576 3023 449578
rect -960 449520 2962 449576
rect 3018 449520 3023 449576
rect -960 449518 3023 449520
rect -960 449428 480 449518
rect 2957 449515 3023 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580441 418298 580507 418301
rect 583520 418298 584960 418388
rect 580441 418296 584960 418298
rect 580441 418240 580446 418296
rect 580502 418240 584960 418296
rect 580441 418238 584960 418240
rect 580441 418235 580507 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3785 397490 3851 397493
rect -960 397488 3851 397490
rect -960 397432 3790 397488
rect 3846 397432 3851 397488
rect -960 397430 3851 397432
rect -960 397340 480 397430
rect 3785 397427 3851 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 578969 378450 579035 378453
rect 583520 378450 584960 378540
rect 578969 378448 584960 378450
rect 578969 378392 578974 378448
rect 579030 378392 584960 378448
rect 578969 378390 584960 378392
rect 578969 378387 579035 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 579981 365122 580047 365125
rect 583520 365122 584960 365212
rect 579981 365120 584960 365122
rect 579981 365064 579986 365120
rect 580042 365064 584960 365120
rect 579981 365062 584960 365064
rect 579981 365059 580047 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2957 345402 3023 345405
rect -960 345400 3023 345402
rect -960 345344 2962 345400
rect 3018 345344 3023 345400
rect -960 345342 3023 345344
rect -960 345252 480 345342
rect 2957 345339 3023 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3233 319290 3299 319293
rect -960 319288 3299 319290
rect -960 319232 3238 319288
rect 3294 319232 3299 319288
rect -960 319230 3299 319232
rect -960 319140 480 319230
rect 3233 319227 3299 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3693 293178 3759 293181
rect -960 293176 3759 293178
rect -960 293120 3698 293176
rect 3754 293120 3759 293176
rect -960 293118 3759 293120
rect -960 293028 480 293118
rect 3693 293115 3759 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 578877 219058 578943 219061
rect 583520 219058 584960 219148
rect 578877 219056 584960 219058
rect 578877 219000 578882 219056
rect 578938 219000 584960 219056
rect 578877 218998 584960 219000
rect 578877 218995 578943 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579889 205730 579955 205733
rect 583520 205730 584960 205820
rect 579889 205728 584960 205730
rect 579889 205672 579894 205728
rect 579950 205672 584960 205728
rect 579889 205670 584960 205672
rect 579889 205667 579955 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 579613 152690 579679 152693
rect 583520 152690 584960 152780
rect 579613 152688 584960 152690
rect 579613 152632 579618 152688
rect 579674 152632 584960 152688
rect 579613 152630 584960 152632
rect 579613 152627 579679 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 580349 139362 580415 139365
rect 583520 139362 584960 139452
rect 580349 139360 584960 139362
rect 580349 139304 580354 139360
rect 580410 139304 584960 139360
rect 580349 139302 584960 139304
rect 580349 139299 580415 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 2773 136778 2839 136781
rect -960 136776 2839 136778
rect -960 136720 2778 136776
rect 2834 136720 2839 136776
rect -960 136718 2839 136720
rect -960 136628 480 136718
rect 2773 136715 2839 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 2957 110666 3023 110669
rect -960 110664 3023 110666
rect -960 110608 2962 110664
rect 3018 110608 3023 110664
rect -960 110606 3023 110608
rect -960 110516 480 110606
rect 2957 110603 3023 110606
rect 580257 99514 580323 99517
rect 583520 99514 584960 99604
rect 580257 99512 584960 99514
rect 580257 99456 580262 99512
rect 580318 99456 584960 99512
rect 580257 99454 584960 99456
rect 580257 99451 580323 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2773 32466 2839 32469
rect -960 32464 2839 32466
rect -960 32408 2778 32464
rect 2834 32408 2839 32464
rect -960 32406 2839 32408
rect -960 32316 480 32406
rect 2773 32403 2839 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 672000 13574 698058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 672000 20414 705242
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 672000 24134 672618
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 672000 27854 676338
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 672000 31574 680058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 672000 38414 686898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 672000 42134 690618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 672000 45854 694338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 672000 49574 698058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 672000 56414 705242
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 672000 60134 672618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 672000 63854 676338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 672000 67574 680058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 672000 74414 686898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 672000 78134 690618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 672000 81854 694338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 672000 85574 698058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 672000 92414 705242
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 672000 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 672000 99854 676338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 672000 103574 680058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 672000 110414 686898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 672000 114134 690618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 672000 117854 694338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 672000 121574 698058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 672000 128414 705242
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 672000 132134 672618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 672000 135854 676338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 672000 139574 680058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 672000 146414 686898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 672000 150134 690618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 672000 153854 694338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 672000 157574 698058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 672000 164414 705242
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 672000 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 672000 171854 676338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 672000 175574 680058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 672000 182414 686898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 672000 186134 690618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 672000 189854 694338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 672000 193574 698058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 672000 200414 705242
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 672000 204134 672618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 672000 207854 676338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 672000 211574 680058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 672000 218414 686898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 672000 222134 690618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 672000 225854 694338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 672000 229574 698058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 672000 236414 705242
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 672000 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 672000 243854 676338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 672000 247574 680058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 672000 254414 686898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 672000 258134 690618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 672000 261854 694338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 672000 265574 698058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 672000 272414 705242
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 672000 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 672000 279854 676338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 672000 283574 680058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 672000 290414 686898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 672000 294134 690618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 672000 297854 694338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 672000 301574 698058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 672000 308414 705242
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 672000 312134 672618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 672000 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 672000 319574 680058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 672000 326414 686898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 672000 330134 690618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 672000 333854 694338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 672000 337574 698058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 672000 344414 705242
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 672000 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 672000 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 672000 355574 680058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 672000 362414 686898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 672000 366134 690618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 672000 369854 694338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 672000 373574 698058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 672000 380414 705242
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 672000 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 672000 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 672000 391574 680058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 672000 398414 686898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 672000 402134 690618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 672000 405854 694338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 672000 409574 698058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 672000 416414 705242
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 672000 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 672000 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 672000 427574 680058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 672000 434414 686898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 672000 438134 690618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 672000 441854 694338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 672000 445574 698058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 672000 452414 705242
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 672000 456134 672618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 672000 459854 676338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 672000 463574 680058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 672000 470414 686898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 672000 474134 690618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 672000 477854 694338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 672000 481574 698058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 672000 488414 705242
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 672000 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 672000 495854 676338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 672000 499574 680058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 672000 506414 686898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 672000 510134 690618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 672000 513854 694338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 672000 517574 698058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 672000 524414 705242
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 672000 528134 672618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 672000 531854 676338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 672000 535574 680058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 672000 542414 686898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 672000 546134 690618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 672000 549854 694338
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 672000 553574 698058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 18208 651454 18528 651486
rect 18208 651218 18250 651454
rect 18486 651218 18528 651454
rect 18208 651134 18528 651218
rect 18208 650898 18250 651134
rect 18486 650898 18528 651134
rect 18208 650866 18528 650898
rect 48928 651454 49248 651486
rect 48928 651218 48970 651454
rect 49206 651218 49248 651454
rect 48928 651134 49248 651218
rect 48928 650898 48970 651134
rect 49206 650898 49248 651134
rect 48928 650866 49248 650898
rect 79648 651454 79968 651486
rect 79648 651218 79690 651454
rect 79926 651218 79968 651454
rect 79648 651134 79968 651218
rect 79648 650898 79690 651134
rect 79926 650898 79968 651134
rect 79648 650866 79968 650898
rect 110368 651454 110688 651486
rect 110368 651218 110410 651454
rect 110646 651218 110688 651454
rect 110368 651134 110688 651218
rect 110368 650898 110410 651134
rect 110646 650898 110688 651134
rect 110368 650866 110688 650898
rect 141088 651454 141408 651486
rect 141088 651218 141130 651454
rect 141366 651218 141408 651454
rect 141088 651134 141408 651218
rect 141088 650898 141130 651134
rect 141366 650898 141408 651134
rect 141088 650866 141408 650898
rect 171808 651454 172128 651486
rect 171808 651218 171850 651454
rect 172086 651218 172128 651454
rect 171808 651134 172128 651218
rect 171808 650898 171850 651134
rect 172086 650898 172128 651134
rect 171808 650866 172128 650898
rect 202528 651454 202848 651486
rect 202528 651218 202570 651454
rect 202806 651218 202848 651454
rect 202528 651134 202848 651218
rect 202528 650898 202570 651134
rect 202806 650898 202848 651134
rect 202528 650866 202848 650898
rect 233248 651454 233568 651486
rect 233248 651218 233290 651454
rect 233526 651218 233568 651454
rect 233248 651134 233568 651218
rect 233248 650898 233290 651134
rect 233526 650898 233568 651134
rect 233248 650866 233568 650898
rect 263968 651454 264288 651486
rect 263968 651218 264010 651454
rect 264246 651218 264288 651454
rect 263968 651134 264288 651218
rect 263968 650898 264010 651134
rect 264246 650898 264288 651134
rect 263968 650866 264288 650898
rect 294688 651454 295008 651486
rect 294688 651218 294730 651454
rect 294966 651218 295008 651454
rect 294688 651134 295008 651218
rect 294688 650898 294730 651134
rect 294966 650898 295008 651134
rect 294688 650866 295008 650898
rect 325408 651454 325728 651486
rect 325408 651218 325450 651454
rect 325686 651218 325728 651454
rect 325408 651134 325728 651218
rect 325408 650898 325450 651134
rect 325686 650898 325728 651134
rect 325408 650866 325728 650898
rect 356128 651454 356448 651486
rect 356128 651218 356170 651454
rect 356406 651218 356448 651454
rect 356128 651134 356448 651218
rect 356128 650898 356170 651134
rect 356406 650898 356448 651134
rect 356128 650866 356448 650898
rect 386848 651454 387168 651486
rect 386848 651218 386890 651454
rect 387126 651218 387168 651454
rect 386848 651134 387168 651218
rect 386848 650898 386890 651134
rect 387126 650898 387168 651134
rect 386848 650866 387168 650898
rect 417568 651454 417888 651486
rect 417568 651218 417610 651454
rect 417846 651218 417888 651454
rect 417568 651134 417888 651218
rect 417568 650898 417610 651134
rect 417846 650898 417888 651134
rect 417568 650866 417888 650898
rect 448288 651454 448608 651486
rect 448288 651218 448330 651454
rect 448566 651218 448608 651454
rect 448288 651134 448608 651218
rect 448288 650898 448330 651134
rect 448566 650898 448608 651134
rect 448288 650866 448608 650898
rect 479008 651454 479328 651486
rect 479008 651218 479050 651454
rect 479286 651218 479328 651454
rect 479008 651134 479328 651218
rect 479008 650898 479050 651134
rect 479286 650898 479328 651134
rect 479008 650866 479328 650898
rect 509728 651454 510048 651486
rect 509728 651218 509770 651454
rect 510006 651218 510048 651454
rect 509728 651134 510048 651218
rect 509728 650898 509770 651134
rect 510006 650898 510048 651134
rect 509728 650866 510048 650898
rect 540448 651454 540768 651486
rect 540448 651218 540490 651454
rect 540726 651218 540768 651454
rect 540448 651134 540768 651218
rect 540448 650898 540490 651134
rect 540726 650898 540768 651134
rect 540448 650866 540768 650898
rect 33568 633454 33888 633486
rect 33568 633218 33610 633454
rect 33846 633218 33888 633454
rect 33568 633134 33888 633218
rect 33568 632898 33610 633134
rect 33846 632898 33888 633134
rect 33568 632866 33888 632898
rect 64288 633454 64608 633486
rect 64288 633218 64330 633454
rect 64566 633218 64608 633454
rect 64288 633134 64608 633218
rect 64288 632898 64330 633134
rect 64566 632898 64608 633134
rect 64288 632866 64608 632898
rect 95008 633454 95328 633486
rect 95008 633218 95050 633454
rect 95286 633218 95328 633454
rect 95008 633134 95328 633218
rect 95008 632898 95050 633134
rect 95286 632898 95328 633134
rect 95008 632866 95328 632898
rect 125728 633454 126048 633486
rect 125728 633218 125770 633454
rect 126006 633218 126048 633454
rect 125728 633134 126048 633218
rect 125728 632898 125770 633134
rect 126006 632898 126048 633134
rect 125728 632866 126048 632898
rect 156448 633454 156768 633486
rect 156448 633218 156490 633454
rect 156726 633218 156768 633454
rect 156448 633134 156768 633218
rect 156448 632898 156490 633134
rect 156726 632898 156768 633134
rect 156448 632866 156768 632898
rect 187168 633454 187488 633486
rect 187168 633218 187210 633454
rect 187446 633218 187488 633454
rect 187168 633134 187488 633218
rect 187168 632898 187210 633134
rect 187446 632898 187488 633134
rect 187168 632866 187488 632898
rect 217888 633454 218208 633486
rect 217888 633218 217930 633454
rect 218166 633218 218208 633454
rect 217888 633134 218208 633218
rect 217888 632898 217930 633134
rect 218166 632898 218208 633134
rect 217888 632866 218208 632898
rect 248608 633454 248928 633486
rect 248608 633218 248650 633454
rect 248886 633218 248928 633454
rect 248608 633134 248928 633218
rect 248608 632898 248650 633134
rect 248886 632898 248928 633134
rect 248608 632866 248928 632898
rect 279328 633454 279648 633486
rect 279328 633218 279370 633454
rect 279606 633218 279648 633454
rect 279328 633134 279648 633218
rect 279328 632898 279370 633134
rect 279606 632898 279648 633134
rect 279328 632866 279648 632898
rect 310048 633454 310368 633486
rect 310048 633218 310090 633454
rect 310326 633218 310368 633454
rect 310048 633134 310368 633218
rect 310048 632898 310090 633134
rect 310326 632898 310368 633134
rect 310048 632866 310368 632898
rect 340768 633454 341088 633486
rect 340768 633218 340810 633454
rect 341046 633218 341088 633454
rect 340768 633134 341088 633218
rect 340768 632898 340810 633134
rect 341046 632898 341088 633134
rect 340768 632866 341088 632898
rect 371488 633454 371808 633486
rect 371488 633218 371530 633454
rect 371766 633218 371808 633454
rect 371488 633134 371808 633218
rect 371488 632898 371530 633134
rect 371766 632898 371808 633134
rect 371488 632866 371808 632898
rect 402208 633454 402528 633486
rect 402208 633218 402250 633454
rect 402486 633218 402528 633454
rect 402208 633134 402528 633218
rect 402208 632898 402250 633134
rect 402486 632898 402528 633134
rect 402208 632866 402528 632898
rect 432928 633454 433248 633486
rect 432928 633218 432970 633454
rect 433206 633218 433248 633454
rect 432928 633134 433248 633218
rect 432928 632898 432970 633134
rect 433206 632898 433248 633134
rect 432928 632866 433248 632898
rect 463648 633454 463968 633486
rect 463648 633218 463690 633454
rect 463926 633218 463968 633454
rect 463648 633134 463968 633218
rect 463648 632898 463690 633134
rect 463926 632898 463968 633134
rect 463648 632866 463968 632898
rect 494368 633454 494688 633486
rect 494368 633218 494410 633454
rect 494646 633218 494688 633454
rect 494368 633134 494688 633218
rect 494368 632898 494410 633134
rect 494646 632898 494688 633134
rect 494368 632866 494688 632898
rect 525088 633454 525408 633486
rect 525088 633218 525130 633454
rect 525366 633218 525408 633454
rect 525088 633134 525408 633218
rect 525088 632898 525130 633134
rect 525366 632898 525408 633134
rect 525088 632866 525408 632898
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 18208 615454 18528 615486
rect 18208 615218 18250 615454
rect 18486 615218 18528 615454
rect 18208 615134 18528 615218
rect 18208 614898 18250 615134
rect 18486 614898 18528 615134
rect 18208 614866 18528 614898
rect 48928 615454 49248 615486
rect 48928 615218 48970 615454
rect 49206 615218 49248 615454
rect 48928 615134 49248 615218
rect 48928 614898 48970 615134
rect 49206 614898 49248 615134
rect 48928 614866 49248 614898
rect 79648 615454 79968 615486
rect 79648 615218 79690 615454
rect 79926 615218 79968 615454
rect 79648 615134 79968 615218
rect 79648 614898 79690 615134
rect 79926 614898 79968 615134
rect 79648 614866 79968 614898
rect 110368 615454 110688 615486
rect 110368 615218 110410 615454
rect 110646 615218 110688 615454
rect 110368 615134 110688 615218
rect 110368 614898 110410 615134
rect 110646 614898 110688 615134
rect 110368 614866 110688 614898
rect 141088 615454 141408 615486
rect 141088 615218 141130 615454
rect 141366 615218 141408 615454
rect 141088 615134 141408 615218
rect 141088 614898 141130 615134
rect 141366 614898 141408 615134
rect 141088 614866 141408 614898
rect 171808 615454 172128 615486
rect 171808 615218 171850 615454
rect 172086 615218 172128 615454
rect 171808 615134 172128 615218
rect 171808 614898 171850 615134
rect 172086 614898 172128 615134
rect 171808 614866 172128 614898
rect 202528 615454 202848 615486
rect 202528 615218 202570 615454
rect 202806 615218 202848 615454
rect 202528 615134 202848 615218
rect 202528 614898 202570 615134
rect 202806 614898 202848 615134
rect 202528 614866 202848 614898
rect 233248 615454 233568 615486
rect 233248 615218 233290 615454
rect 233526 615218 233568 615454
rect 233248 615134 233568 615218
rect 233248 614898 233290 615134
rect 233526 614898 233568 615134
rect 233248 614866 233568 614898
rect 263968 615454 264288 615486
rect 263968 615218 264010 615454
rect 264246 615218 264288 615454
rect 263968 615134 264288 615218
rect 263968 614898 264010 615134
rect 264246 614898 264288 615134
rect 263968 614866 264288 614898
rect 294688 615454 295008 615486
rect 294688 615218 294730 615454
rect 294966 615218 295008 615454
rect 294688 615134 295008 615218
rect 294688 614898 294730 615134
rect 294966 614898 295008 615134
rect 294688 614866 295008 614898
rect 325408 615454 325728 615486
rect 325408 615218 325450 615454
rect 325686 615218 325728 615454
rect 325408 615134 325728 615218
rect 325408 614898 325450 615134
rect 325686 614898 325728 615134
rect 325408 614866 325728 614898
rect 356128 615454 356448 615486
rect 356128 615218 356170 615454
rect 356406 615218 356448 615454
rect 356128 615134 356448 615218
rect 356128 614898 356170 615134
rect 356406 614898 356448 615134
rect 356128 614866 356448 614898
rect 386848 615454 387168 615486
rect 386848 615218 386890 615454
rect 387126 615218 387168 615454
rect 386848 615134 387168 615218
rect 386848 614898 386890 615134
rect 387126 614898 387168 615134
rect 386848 614866 387168 614898
rect 417568 615454 417888 615486
rect 417568 615218 417610 615454
rect 417846 615218 417888 615454
rect 417568 615134 417888 615218
rect 417568 614898 417610 615134
rect 417846 614898 417888 615134
rect 417568 614866 417888 614898
rect 448288 615454 448608 615486
rect 448288 615218 448330 615454
rect 448566 615218 448608 615454
rect 448288 615134 448608 615218
rect 448288 614898 448330 615134
rect 448566 614898 448608 615134
rect 448288 614866 448608 614898
rect 479008 615454 479328 615486
rect 479008 615218 479050 615454
rect 479286 615218 479328 615454
rect 479008 615134 479328 615218
rect 479008 614898 479050 615134
rect 479286 614898 479328 615134
rect 479008 614866 479328 614898
rect 509728 615454 510048 615486
rect 509728 615218 509770 615454
rect 510006 615218 510048 615454
rect 509728 615134 510048 615218
rect 509728 614898 509770 615134
rect 510006 614898 510048 615134
rect 509728 614866 510048 614898
rect 540448 615454 540768 615486
rect 540448 615218 540490 615454
rect 540726 615218 540768 615454
rect 540448 615134 540768 615218
rect 540448 614898 540490 615134
rect 540726 614898 540768 615134
rect 540448 614866 540768 614898
rect 33568 597454 33888 597486
rect 33568 597218 33610 597454
rect 33846 597218 33888 597454
rect 33568 597134 33888 597218
rect 33568 596898 33610 597134
rect 33846 596898 33888 597134
rect 33568 596866 33888 596898
rect 64288 597454 64608 597486
rect 64288 597218 64330 597454
rect 64566 597218 64608 597454
rect 64288 597134 64608 597218
rect 64288 596898 64330 597134
rect 64566 596898 64608 597134
rect 64288 596866 64608 596898
rect 95008 597454 95328 597486
rect 95008 597218 95050 597454
rect 95286 597218 95328 597454
rect 95008 597134 95328 597218
rect 95008 596898 95050 597134
rect 95286 596898 95328 597134
rect 95008 596866 95328 596898
rect 125728 597454 126048 597486
rect 125728 597218 125770 597454
rect 126006 597218 126048 597454
rect 125728 597134 126048 597218
rect 125728 596898 125770 597134
rect 126006 596898 126048 597134
rect 125728 596866 126048 596898
rect 156448 597454 156768 597486
rect 156448 597218 156490 597454
rect 156726 597218 156768 597454
rect 156448 597134 156768 597218
rect 156448 596898 156490 597134
rect 156726 596898 156768 597134
rect 156448 596866 156768 596898
rect 187168 597454 187488 597486
rect 187168 597218 187210 597454
rect 187446 597218 187488 597454
rect 187168 597134 187488 597218
rect 187168 596898 187210 597134
rect 187446 596898 187488 597134
rect 187168 596866 187488 596898
rect 217888 597454 218208 597486
rect 217888 597218 217930 597454
rect 218166 597218 218208 597454
rect 217888 597134 218208 597218
rect 217888 596898 217930 597134
rect 218166 596898 218208 597134
rect 217888 596866 218208 596898
rect 248608 597454 248928 597486
rect 248608 597218 248650 597454
rect 248886 597218 248928 597454
rect 248608 597134 248928 597218
rect 248608 596898 248650 597134
rect 248886 596898 248928 597134
rect 248608 596866 248928 596898
rect 279328 597454 279648 597486
rect 279328 597218 279370 597454
rect 279606 597218 279648 597454
rect 279328 597134 279648 597218
rect 279328 596898 279370 597134
rect 279606 596898 279648 597134
rect 279328 596866 279648 596898
rect 310048 597454 310368 597486
rect 310048 597218 310090 597454
rect 310326 597218 310368 597454
rect 310048 597134 310368 597218
rect 310048 596898 310090 597134
rect 310326 596898 310368 597134
rect 310048 596866 310368 596898
rect 340768 597454 341088 597486
rect 340768 597218 340810 597454
rect 341046 597218 341088 597454
rect 340768 597134 341088 597218
rect 340768 596898 340810 597134
rect 341046 596898 341088 597134
rect 340768 596866 341088 596898
rect 371488 597454 371808 597486
rect 371488 597218 371530 597454
rect 371766 597218 371808 597454
rect 371488 597134 371808 597218
rect 371488 596898 371530 597134
rect 371766 596898 371808 597134
rect 371488 596866 371808 596898
rect 402208 597454 402528 597486
rect 402208 597218 402250 597454
rect 402486 597218 402528 597454
rect 402208 597134 402528 597218
rect 402208 596898 402250 597134
rect 402486 596898 402528 597134
rect 402208 596866 402528 596898
rect 432928 597454 433248 597486
rect 432928 597218 432970 597454
rect 433206 597218 433248 597454
rect 432928 597134 433248 597218
rect 432928 596898 432970 597134
rect 433206 596898 433248 597134
rect 432928 596866 433248 596898
rect 463648 597454 463968 597486
rect 463648 597218 463690 597454
rect 463926 597218 463968 597454
rect 463648 597134 463968 597218
rect 463648 596898 463690 597134
rect 463926 596898 463968 597134
rect 463648 596866 463968 596898
rect 494368 597454 494688 597486
rect 494368 597218 494410 597454
rect 494646 597218 494688 597454
rect 494368 597134 494688 597218
rect 494368 596898 494410 597134
rect 494646 596898 494688 597134
rect 494368 596866 494688 596898
rect 525088 597454 525408 597486
rect 525088 597218 525130 597454
rect 525366 597218 525408 597454
rect 525088 597134 525408 597218
rect 525088 596898 525130 597134
rect 525366 596898 525408 597134
rect 525088 596866 525408 596898
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 18208 579454 18528 579486
rect 18208 579218 18250 579454
rect 18486 579218 18528 579454
rect 18208 579134 18528 579218
rect 18208 578898 18250 579134
rect 18486 578898 18528 579134
rect 18208 578866 18528 578898
rect 48928 579454 49248 579486
rect 48928 579218 48970 579454
rect 49206 579218 49248 579454
rect 48928 579134 49248 579218
rect 48928 578898 48970 579134
rect 49206 578898 49248 579134
rect 48928 578866 49248 578898
rect 79648 579454 79968 579486
rect 79648 579218 79690 579454
rect 79926 579218 79968 579454
rect 79648 579134 79968 579218
rect 79648 578898 79690 579134
rect 79926 578898 79968 579134
rect 79648 578866 79968 578898
rect 110368 579454 110688 579486
rect 110368 579218 110410 579454
rect 110646 579218 110688 579454
rect 110368 579134 110688 579218
rect 110368 578898 110410 579134
rect 110646 578898 110688 579134
rect 110368 578866 110688 578898
rect 141088 579454 141408 579486
rect 141088 579218 141130 579454
rect 141366 579218 141408 579454
rect 141088 579134 141408 579218
rect 141088 578898 141130 579134
rect 141366 578898 141408 579134
rect 141088 578866 141408 578898
rect 171808 579454 172128 579486
rect 171808 579218 171850 579454
rect 172086 579218 172128 579454
rect 171808 579134 172128 579218
rect 171808 578898 171850 579134
rect 172086 578898 172128 579134
rect 171808 578866 172128 578898
rect 202528 579454 202848 579486
rect 202528 579218 202570 579454
rect 202806 579218 202848 579454
rect 202528 579134 202848 579218
rect 202528 578898 202570 579134
rect 202806 578898 202848 579134
rect 202528 578866 202848 578898
rect 233248 579454 233568 579486
rect 233248 579218 233290 579454
rect 233526 579218 233568 579454
rect 233248 579134 233568 579218
rect 233248 578898 233290 579134
rect 233526 578898 233568 579134
rect 233248 578866 233568 578898
rect 263968 579454 264288 579486
rect 263968 579218 264010 579454
rect 264246 579218 264288 579454
rect 263968 579134 264288 579218
rect 263968 578898 264010 579134
rect 264246 578898 264288 579134
rect 263968 578866 264288 578898
rect 294688 579454 295008 579486
rect 294688 579218 294730 579454
rect 294966 579218 295008 579454
rect 294688 579134 295008 579218
rect 294688 578898 294730 579134
rect 294966 578898 295008 579134
rect 294688 578866 295008 578898
rect 325408 579454 325728 579486
rect 325408 579218 325450 579454
rect 325686 579218 325728 579454
rect 325408 579134 325728 579218
rect 325408 578898 325450 579134
rect 325686 578898 325728 579134
rect 325408 578866 325728 578898
rect 356128 579454 356448 579486
rect 356128 579218 356170 579454
rect 356406 579218 356448 579454
rect 356128 579134 356448 579218
rect 356128 578898 356170 579134
rect 356406 578898 356448 579134
rect 356128 578866 356448 578898
rect 386848 579454 387168 579486
rect 386848 579218 386890 579454
rect 387126 579218 387168 579454
rect 386848 579134 387168 579218
rect 386848 578898 386890 579134
rect 387126 578898 387168 579134
rect 386848 578866 387168 578898
rect 417568 579454 417888 579486
rect 417568 579218 417610 579454
rect 417846 579218 417888 579454
rect 417568 579134 417888 579218
rect 417568 578898 417610 579134
rect 417846 578898 417888 579134
rect 417568 578866 417888 578898
rect 448288 579454 448608 579486
rect 448288 579218 448330 579454
rect 448566 579218 448608 579454
rect 448288 579134 448608 579218
rect 448288 578898 448330 579134
rect 448566 578898 448608 579134
rect 448288 578866 448608 578898
rect 479008 579454 479328 579486
rect 479008 579218 479050 579454
rect 479286 579218 479328 579454
rect 479008 579134 479328 579218
rect 479008 578898 479050 579134
rect 479286 578898 479328 579134
rect 479008 578866 479328 578898
rect 509728 579454 510048 579486
rect 509728 579218 509770 579454
rect 510006 579218 510048 579454
rect 509728 579134 510048 579218
rect 509728 578898 509770 579134
rect 510006 578898 510048 579134
rect 509728 578866 510048 578898
rect 540448 579454 540768 579486
rect 540448 579218 540490 579454
rect 540726 579218 540768 579454
rect 540448 579134 540768 579218
rect 540448 578898 540490 579134
rect 540726 578898 540768 579134
rect 540448 578866 540768 578898
rect 33568 561454 33888 561486
rect 33568 561218 33610 561454
rect 33846 561218 33888 561454
rect 33568 561134 33888 561218
rect 33568 560898 33610 561134
rect 33846 560898 33888 561134
rect 33568 560866 33888 560898
rect 64288 561454 64608 561486
rect 64288 561218 64330 561454
rect 64566 561218 64608 561454
rect 64288 561134 64608 561218
rect 64288 560898 64330 561134
rect 64566 560898 64608 561134
rect 64288 560866 64608 560898
rect 95008 561454 95328 561486
rect 95008 561218 95050 561454
rect 95286 561218 95328 561454
rect 95008 561134 95328 561218
rect 95008 560898 95050 561134
rect 95286 560898 95328 561134
rect 95008 560866 95328 560898
rect 125728 561454 126048 561486
rect 125728 561218 125770 561454
rect 126006 561218 126048 561454
rect 125728 561134 126048 561218
rect 125728 560898 125770 561134
rect 126006 560898 126048 561134
rect 125728 560866 126048 560898
rect 156448 561454 156768 561486
rect 156448 561218 156490 561454
rect 156726 561218 156768 561454
rect 156448 561134 156768 561218
rect 156448 560898 156490 561134
rect 156726 560898 156768 561134
rect 156448 560866 156768 560898
rect 187168 561454 187488 561486
rect 187168 561218 187210 561454
rect 187446 561218 187488 561454
rect 187168 561134 187488 561218
rect 187168 560898 187210 561134
rect 187446 560898 187488 561134
rect 187168 560866 187488 560898
rect 217888 561454 218208 561486
rect 217888 561218 217930 561454
rect 218166 561218 218208 561454
rect 217888 561134 218208 561218
rect 217888 560898 217930 561134
rect 218166 560898 218208 561134
rect 217888 560866 218208 560898
rect 248608 561454 248928 561486
rect 248608 561218 248650 561454
rect 248886 561218 248928 561454
rect 248608 561134 248928 561218
rect 248608 560898 248650 561134
rect 248886 560898 248928 561134
rect 248608 560866 248928 560898
rect 279328 561454 279648 561486
rect 279328 561218 279370 561454
rect 279606 561218 279648 561454
rect 279328 561134 279648 561218
rect 279328 560898 279370 561134
rect 279606 560898 279648 561134
rect 279328 560866 279648 560898
rect 310048 561454 310368 561486
rect 310048 561218 310090 561454
rect 310326 561218 310368 561454
rect 310048 561134 310368 561218
rect 310048 560898 310090 561134
rect 310326 560898 310368 561134
rect 310048 560866 310368 560898
rect 340768 561454 341088 561486
rect 340768 561218 340810 561454
rect 341046 561218 341088 561454
rect 340768 561134 341088 561218
rect 340768 560898 340810 561134
rect 341046 560898 341088 561134
rect 340768 560866 341088 560898
rect 371488 561454 371808 561486
rect 371488 561218 371530 561454
rect 371766 561218 371808 561454
rect 371488 561134 371808 561218
rect 371488 560898 371530 561134
rect 371766 560898 371808 561134
rect 371488 560866 371808 560898
rect 402208 561454 402528 561486
rect 402208 561218 402250 561454
rect 402486 561218 402528 561454
rect 402208 561134 402528 561218
rect 402208 560898 402250 561134
rect 402486 560898 402528 561134
rect 402208 560866 402528 560898
rect 432928 561454 433248 561486
rect 432928 561218 432970 561454
rect 433206 561218 433248 561454
rect 432928 561134 433248 561218
rect 432928 560898 432970 561134
rect 433206 560898 433248 561134
rect 432928 560866 433248 560898
rect 463648 561454 463968 561486
rect 463648 561218 463690 561454
rect 463926 561218 463968 561454
rect 463648 561134 463968 561218
rect 463648 560898 463690 561134
rect 463926 560898 463968 561134
rect 463648 560866 463968 560898
rect 494368 561454 494688 561486
rect 494368 561218 494410 561454
rect 494646 561218 494688 561454
rect 494368 561134 494688 561218
rect 494368 560898 494410 561134
rect 494646 560898 494688 561134
rect 494368 560866 494688 560898
rect 525088 561454 525408 561486
rect 525088 561218 525130 561454
rect 525366 561218 525408 561454
rect 525088 561134 525408 561218
rect 525088 560898 525130 561134
rect 525366 560898 525408 561134
rect 525088 560866 525408 560898
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 18208 543454 18528 543486
rect 18208 543218 18250 543454
rect 18486 543218 18528 543454
rect 18208 543134 18528 543218
rect 18208 542898 18250 543134
rect 18486 542898 18528 543134
rect 18208 542866 18528 542898
rect 48928 543454 49248 543486
rect 48928 543218 48970 543454
rect 49206 543218 49248 543454
rect 48928 543134 49248 543218
rect 48928 542898 48970 543134
rect 49206 542898 49248 543134
rect 48928 542866 49248 542898
rect 79648 543454 79968 543486
rect 79648 543218 79690 543454
rect 79926 543218 79968 543454
rect 79648 543134 79968 543218
rect 79648 542898 79690 543134
rect 79926 542898 79968 543134
rect 79648 542866 79968 542898
rect 110368 543454 110688 543486
rect 110368 543218 110410 543454
rect 110646 543218 110688 543454
rect 110368 543134 110688 543218
rect 110368 542898 110410 543134
rect 110646 542898 110688 543134
rect 110368 542866 110688 542898
rect 141088 543454 141408 543486
rect 141088 543218 141130 543454
rect 141366 543218 141408 543454
rect 141088 543134 141408 543218
rect 141088 542898 141130 543134
rect 141366 542898 141408 543134
rect 141088 542866 141408 542898
rect 171808 543454 172128 543486
rect 171808 543218 171850 543454
rect 172086 543218 172128 543454
rect 171808 543134 172128 543218
rect 171808 542898 171850 543134
rect 172086 542898 172128 543134
rect 171808 542866 172128 542898
rect 202528 543454 202848 543486
rect 202528 543218 202570 543454
rect 202806 543218 202848 543454
rect 202528 543134 202848 543218
rect 202528 542898 202570 543134
rect 202806 542898 202848 543134
rect 202528 542866 202848 542898
rect 233248 543454 233568 543486
rect 233248 543218 233290 543454
rect 233526 543218 233568 543454
rect 233248 543134 233568 543218
rect 233248 542898 233290 543134
rect 233526 542898 233568 543134
rect 233248 542866 233568 542898
rect 263968 543454 264288 543486
rect 263968 543218 264010 543454
rect 264246 543218 264288 543454
rect 263968 543134 264288 543218
rect 263968 542898 264010 543134
rect 264246 542898 264288 543134
rect 263968 542866 264288 542898
rect 294688 543454 295008 543486
rect 294688 543218 294730 543454
rect 294966 543218 295008 543454
rect 294688 543134 295008 543218
rect 294688 542898 294730 543134
rect 294966 542898 295008 543134
rect 294688 542866 295008 542898
rect 325408 543454 325728 543486
rect 325408 543218 325450 543454
rect 325686 543218 325728 543454
rect 325408 543134 325728 543218
rect 325408 542898 325450 543134
rect 325686 542898 325728 543134
rect 325408 542866 325728 542898
rect 356128 543454 356448 543486
rect 356128 543218 356170 543454
rect 356406 543218 356448 543454
rect 356128 543134 356448 543218
rect 356128 542898 356170 543134
rect 356406 542898 356448 543134
rect 356128 542866 356448 542898
rect 386848 543454 387168 543486
rect 386848 543218 386890 543454
rect 387126 543218 387168 543454
rect 386848 543134 387168 543218
rect 386848 542898 386890 543134
rect 387126 542898 387168 543134
rect 386848 542866 387168 542898
rect 417568 543454 417888 543486
rect 417568 543218 417610 543454
rect 417846 543218 417888 543454
rect 417568 543134 417888 543218
rect 417568 542898 417610 543134
rect 417846 542898 417888 543134
rect 417568 542866 417888 542898
rect 448288 543454 448608 543486
rect 448288 543218 448330 543454
rect 448566 543218 448608 543454
rect 448288 543134 448608 543218
rect 448288 542898 448330 543134
rect 448566 542898 448608 543134
rect 448288 542866 448608 542898
rect 479008 543454 479328 543486
rect 479008 543218 479050 543454
rect 479286 543218 479328 543454
rect 479008 543134 479328 543218
rect 479008 542898 479050 543134
rect 479286 542898 479328 543134
rect 479008 542866 479328 542898
rect 509728 543454 510048 543486
rect 509728 543218 509770 543454
rect 510006 543218 510048 543454
rect 509728 543134 510048 543218
rect 509728 542898 509770 543134
rect 510006 542898 510048 543134
rect 509728 542866 510048 542898
rect 540448 543454 540768 543486
rect 540448 543218 540490 543454
rect 540726 543218 540768 543454
rect 540448 543134 540768 543218
rect 540448 542898 540490 543134
rect 540726 542898 540768 543134
rect 540448 542866 540768 542898
rect 33568 525454 33888 525486
rect 33568 525218 33610 525454
rect 33846 525218 33888 525454
rect 33568 525134 33888 525218
rect 33568 524898 33610 525134
rect 33846 524898 33888 525134
rect 33568 524866 33888 524898
rect 64288 525454 64608 525486
rect 64288 525218 64330 525454
rect 64566 525218 64608 525454
rect 64288 525134 64608 525218
rect 64288 524898 64330 525134
rect 64566 524898 64608 525134
rect 64288 524866 64608 524898
rect 95008 525454 95328 525486
rect 95008 525218 95050 525454
rect 95286 525218 95328 525454
rect 95008 525134 95328 525218
rect 95008 524898 95050 525134
rect 95286 524898 95328 525134
rect 95008 524866 95328 524898
rect 125728 525454 126048 525486
rect 125728 525218 125770 525454
rect 126006 525218 126048 525454
rect 125728 525134 126048 525218
rect 125728 524898 125770 525134
rect 126006 524898 126048 525134
rect 125728 524866 126048 524898
rect 156448 525454 156768 525486
rect 156448 525218 156490 525454
rect 156726 525218 156768 525454
rect 156448 525134 156768 525218
rect 156448 524898 156490 525134
rect 156726 524898 156768 525134
rect 156448 524866 156768 524898
rect 187168 525454 187488 525486
rect 187168 525218 187210 525454
rect 187446 525218 187488 525454
rect 187168 525134 187488 525218
rect 187168 524898 187210 525134
rect 187446 524898 187488 525134
rect 187168 524866 187488 524898
rect 217888 525454 218208 525486
rect 217888 525218 217930 525454
rect 218166 525218 218208 525454
rect 217888 525134 218208 525218
rect 217888 524898 217930 525134
rect 218166 524898 218208 525134
rect 217888 524866 218208 524898
rect 248608 525454 248928 525486
rect 248608 525218 248650 525454
rect 248886 525218 248928 525454
rect 248608 525134 248928 525218
rect 248608 524898 248650 525134
rect 248886 524898 248928 525134
rect 248608 524866 248928 524898
rect 279328 525454 279648 525486
rect 279328 525218 279370 525454
rect 279606 525218 279648 525454
rect 279328 525134 279648 525218
rect 279328 524898 279370 525134
rect 279606 524898 279648 525134
rect 279328 524866 279648 524898
rect 310048 525454 310368 525486
rect 310048 525218 310090 525454
rect 310326 525218 310368 525454
rect 310048 525134 310368 525218
rect 310048 524898 310090 525134
rect 310326 524898 310368 525134
rect 310048 524866 310368 524898
rect 340768 525454 341088 525486
rect 340768 525218 340810 525454
rect 341046 525218 341088 525454
rect 340768 525134 341088 525218
rect 340768 524898 340810 525134
rect 341046 524898 341088 525134
rect 340768 524866 341088 524898
rect 371488 525454 371808 525486
rect 371488 525218 371530 525454
rect 371766 525218 371808 525454
rect 371488 525134 371808 525218
rect 371488 524898 371530 525134
rect 371766 524898 371808 525134
rect 371488 524866 371808 524898
rect 402208 525454 402528 525486
rect 402208 525218 402250 525454
rect 402486 525218 402528 525454
rect 402208 525134 402528 525218
rect 402208 524898 402250 525134
rect 402486 524898 402528 525134
rect 402208 524866 402528 524898
rect 432928 525454 433248 525486
rect 432928 525218 432970 525454
rect 433206 525218 433248 525454
rect 432928 525134 433248 525218
rect 432928 524898 432970 525134
rect 433206 524898 433248 525134
rect 432928 524866 433248 524898
rect 463648 525454 463968 525486
rect 463648 525218 463690 525454
rect 463926 525218 463968 525454
rect 463648 525134 463968 525218
rect 463648 524898 463690 525134
rect 463926 524898 463968 525134
rect 463648 524866 463968 524898
rect 494368 525454 494688 525486
rect 494368 525218 494410 525454
rect 494646 525218 494688 525454
rect 494368 525134 494688 525218
rect 494368 524898 494410 525134
rect 494646 524898 494688 525134
rect 494368 524866 494688 524898
rect 525088 525454 525408 525486
rect 525088 525218 525130 525454
rect 525366 525218 525408 525454
rect 525088 525134 525408 525218
rect 525088 524898 525130 525134
rect 525366 524898 525408 525134
rect 525088 524866 525408 524898
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 18208 507454 18528 507486
rect 18208 507218 18250 507454
rect 18486 507218 18528 507454
rect 18208 507134 18528 507218
rect 18208 506898 18250 507134
rect 18486 506898 18528 507134
rect 18208 506866 18528 506898
rect 48928 507454 49248 507486
rect 48928 507218 48970 507454
rect 49206 507218 49248 507454
rect 48928 507134 49248 507218
rect 48928 506898 48970 507134
rect 49206 506898 49248 507134
rect 48928 506866 49248 506898
rect 79648 507454 79968 507486
rect 79648 507218 79690 507454
rect 79926 507218 79968 507454
rect 79648 507134 79968 507218
rect 79648 506898 79690 507134
rect 79926 506898 79968 507134
rect 79648 506866 79968 506898
rect 110368 507454 110688 507486
rect 110368 507218 110410 507454
rect 110646 507218 110688 507454
rect 110368 507134 110688 507218
rect 110368 506898 110410 507134
rect 110646 506898 110688 507134
rect 110368 506866 110688 506898
rect 141088 507454 141408 507486
rect 141088 507218 141130 507454
rect 141366 507218 141408 507454
rect 141088 507134 141408 507218
rect 141088 506898 141130 507134
rect 141366 506898 141408 507134
rect 141088 506866 141408 506898
rect 171808 507454 172128 507486
rect 171808 507218 171850 507454
rect 172086 507218 172128 507454
rect 171808 507134 172128 507218
rect 171808 506898 171850 507134
rect 172086 506898 172128 507134
rect 171808 506866 172128 506898
rect 202528 507454 202848 507486
rect 202528 507218 202570 507454
rect 202806 507218 202848 507454
rect 202528 507134 202848 507218
rect 202528 506898 202570 507134
rect 202806 506898 202848 507134
rect 202528 506866 202848 506898
rect 233248 507454 233568 507486
rect 233248 507218 233290 507454
rect 233526 507218 233568 507454
rect 233248 507134 233568 507218
rect 233248 506898 233290 507134
rect 233526 506898 233568 507134
rect 233248 506866 233568 506898
rect 263968 507454 264288 507486
rect 263968 507218 264010 507454
rect 264246 507218 264288 507454
rect 263968 507134 264288 507218
rect 263968 506898 264010 507134
rect 264246 506898 264288 507134
rect 263968 506866 264288 506898
rect 294688 507454 295008 507486
rect 294688 507218 294730 507454
rect 294966 507218 295008 507454
rect 294688 507134 295008 507218
rect 294688 506898 294730 507134
rect 294966 506898 295008 507134
rect 294688 506866 295008 506898
rect 325408 507454 325728 507486
rect 325408 507218 325450 507454
rect 325686 507218 325728 507454
rect 325408 507134 325728 507218
rect 325408 506898 325450 507134
rect 325686 506898 325728 507134
rect 325408 506866 325728 506898
rect 356128 507454 356448 507486
rect 356128 507218 356170 507454
rect 356406 507218 356448 507454
rect 356128 507134 356448 507218
rect 356128 506898 356170 507134
rect 356406 506898 356448 507134
rect 356128 506866 356448 506898
rect 386848 507454 387168 507486
rect 386848 507218 386890 507454
rect 387126 507218 387168 507454
rect 386848 507134 387168 507218
rect 386848 506898 386890 507134
rect 387126 506898 387168 507134
rect 386848 506866 387168 506898
rect 417568 507454 417888 507486
rect 417568 507218 417610 507454
rect 417846 507218 417888 507454
rect 417568 507134 417888 507218
rect 417568 506898 417610 507134
rect 417846 506898 417888 507134
rect 417568 506866 417888 506898
rect 448288 507454 448608 507486
rect 448288 507218 448330 507454
rect 448566 507218 448608 507454
rect 448288 507134 448608 507218
rect 448288 506898 448330 507134
rect 448566 506898 448608 507134
rect 448288 506866 448608 506898
rect 479008 507454 479328 507486
rect 479008 507218 479050 507454
rect 479286 507218 479328 507454
rect 479008 507134 479328 507218
rect 479008 506898 479050 507134
rect 479286 506898 479328 507134
rect 479008 506866 479328 506898
rect 509728 507454 510048 507486
rect 509728 507218 509770 507454
rect 510006 507218 510048 507454
rect 509728 507134 510048 507218
rect 509728 506898 509770 507134
rect 510006 506898 510048 507134
rect 509728 506866 510048 506898
rect 540448 507454 540768 507486
rect 540448 507218 540490 507454
rect 540726 507218 540768 507454
rect 540448 507134 540768 507218
rect 540448 506898 540490 507134
rect 540726 506898 540768 507134
rect 540448 506866 540768 506898
rect 33568 489454 33888 489486
rect 33568 489218 33610 489454
rect 33846 489218 33888 489454
rect 33568 489134 33888 489218
rect 33568 488898 33610 489134
rect 33846 488898 33888 489134
rect 33568 488866 33888 488898
rect 64288 489454 64608 489486
rect 64288 489218 64330 489454
rect 64566 489218 64608 489454
rect 64288 489134 64608 489218
rect 64288 488898 64330 489134
rect 64566 488898 64608 489134
rect 64288 488866 64608 488898
rect 95008 489454 95328 489486
rect 95008 489218 95050 489454
rect 95286 489218 95328 489454
rect 95008 489134 95328 489218
rect 95008 488898 95050 489134
rect 95286 488898 95328 489134
rect 95008 488866 95328 488898
rect 125728 489454 126048 489486
rect 125728 489218 125770 489454
rect 126006 489218 126048 489454
rect 125728 489134 126048 489218
rect 125728 488898 125770 489134
rect 126006 488898 126048 489134
rect 125728 488866 126048 488898
rect 156448 489454 156768 489486
rect 156448 489218 156490 489454
rect 156726 489218 156768 489454
rect 156448 489134 156768 489218
rect 156448 488898 156490 489134
rect 156726 488898 156768 489134
rect 156448 488866 156768 488898
rect 187168 489454 187488 489486
rect 187168 489218 187210 489454
rect 187446 489218 187488 489454
rect 187168 489134 187488 489218
rect 187168 488898 187210 489134
rect 187446 488898 187488 489134
rect 187168 488866 187488 488898
rect 217888 489454 218208 489486
rect 217888 489218 217930 489454
rect 218166 489218 218208 489454
rect 217888 489134 218208 489218
rect 217888 488898 217930 489134
rect 218166 488898 218208 489134
rect 217888 488866 218208 488898
rect 248608 489454 248928 489486
rect 248608 489218 248650 489454
rect 248886 489218 248928 489454
rect 248608 489134 248928 489218
rect 248608 488898 248650 489134
rect 248886 488898 248928 489134
rect 248608 488866 248928 488898
rect 279328 489454 279648 489486
rect 279328 489218 279370 489454
rect 279606 489218 279648 489454
rect 279328 489134 279648 489218
rect 279328 488898 279370 489134
rect 279606 488898 279648 489134
rect 279328 488866 279648 488898
rect 310048 489454 310368 489486
rect 310048 489218 310090 489454
rect 310326 489218 310368 489454
rect 310048 489134 310368 489218
rect 310048 488898 310090 489134
rect 310326 488898 310368 489134
rect 310048 488866 310368 488898
rect 340768 489454 341088 489486
rect 340768 489218 340810 489454
rect 341046 489218 341088 489454
rect 340768 489134 341088 489218
rect 340768 488898 340810 489134
rect 341046 488898 341088 489134
rect 340768 488866 341088 488898
rect 371488 489454 371808 489486
rect 371488 489218 371530 489454
rect 371766 489218 371808 489454
rect 371488 489134 371808 489218
rect 371488 488898 371530 489134
rect 371766 488898 371808 489134
rect 371488 488866 371808 488898
rect 402208 489454 402528 489486
rect 402208 489218 402250 489454
rect 402486 489218 402528 489454
rect 402208 489134 402528 489218
rect 402208 488898 402250 489134
rect 402486 488898 402528 489134
rect 402208 488866 402528 488898
rect 432928 489454 433248 489486
rect 432928 489218 432970 489454
rect 433206 489218 433248 489454
rect 432928 489134 433248 489218
rect 432928 488898 432970 489134
rect 433206 488898 433248 489134
rect 432928 488866 433248 488898
rect 463648 489454 463968 489486
rect 463648 489218 463690 489454
rect 463926 489218 463968 489454
rect 463648 489134 463968 489218
rect 463648 488898 463690 489134
rect 463926 488898 463968 489134
rect 463648 488866 463968 488898
rect 494368 489454 494688 489486
rect 494368 489218 494410 489454
rect 494646 489218 494688 489454
rect 494368 489134 494688 489218
rect 494368 488898 494410 489134
rect 494646 488898 494688 489134
rect 494368 488866 494688 488898
rect 525088 489454 525408 489486
rect 525088 489218 525130 489454
rect 525366 489218 525408 489454
rect 525088 489134 525408 489218
rect 525088 488898 525130 489134
rect 525366 488898 525408 489134
rect 525088 488866 525408 488898
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 18208 471454 18528 471486
rect 18208 471218 18250 471454
rect 18486 471218 18528 471454
rect 18208 471134 18528 471218
rect 18208 470898 18250 471134
rect 18486 470898 18528 471134
rect 18208 470866 18528 470898
rect 48928 471454 49248 471486
rect 48928 471218 48970 471454
rect 49206 471218 49248 471454
rect 48928 471134 49248 471218
rect 48928 470898 48970 471134
rect 49206 470898 49248 471134
rect 48928 470866 49248 470898
rect 79648 471454 79968 471486
rect 79648 471218 79690 471454
rect 79926 471218 79968 471454
rect 79648 471134 79968 471218
rect 79648 470898 79690 471134
rect 79926 470898 79968 471134
rect 79648 470866 79968 470898
rect 110368 471454 110688 471486
rect 110368 471218 110410 471454
rect 110646 471218 110688 471454
rect 110368 471134 110688 471218
rect 110368 470898 110410 471134
rect 110646 470898 110688 471134
rect 110368 470866 110688 470898
rect 141088 471454 141408 471486
rect 141088 471218 141130 471454
rect 141366 471218 141408 471454
rect 141088 471134 141408 471218
rect 141088 470898 141130 471134
rect 141366 470898 141408 471134
rect 141088 470866 141408 470898
rect 171808 471454 172128 471486
rect 171808 471218 171850 471454
rect 172086 471218 172128 471454
rect 171808 471134 172128 471218
rect 171808 470898 171850 471134
rect 172086 470898 172128 471134
rect 171808 470866 172128 470898
rect 202528 471454 202848 471486
rect 202528 471218 202570 471454
rect 202806 471218 202848 471454
rect 202528 471134 202848 471218
rect 202528 470898 202570 471134
rect 202806 470898 202848 471134
rect 202528 470866 202848 470898
rect 233248 471454 233568 471486
rect 233248 471218 233290 471454
rect 233526 471218 233568 471454
rect 233248 471134 233568 471218
rect 233248 470898 233290 471134
rect 233526 470898 233568 471134
rect 233248 470866 233568 470898
rect 263968 471454 264288 471486
rect 263968 471218 264010 471454
rect 264246 471218 264288 471454
rect 263968 471134 264288 471218
rect 263968 470898 264010 471134
rect 264246 470898 264288 471134
rect 263968 470866 264288 470898
rect 294688 471454 295008 471486
rect 294688 471218 294730 471454
rect 294966 471218 295008 471454
rect 294688 471134 295008 471218
rect 294688 470898 294730 471134
rect 294966 470898 295008 471134
rect 294688 470866 295008 470898
rect 325408 471454 325728 471486
rect 325408 471218 325450 471454
rect 325686 471218 325728 471454
rect 325408 471134 325728 471218
rect 325408 470898 325450 471134
rect 325686 470898 325728 471134
rect 325408 470866 325728 470898
rect 356128 471454 356448 471486
rect 356128 471218 356170 471454
rect 356406 471218 356448 471454
rect 356128 471134 356448 471218
rect 356128 470898 356170 471134
rect 356406 470898 356448 471134
rect 356128 470866 356448 470898
rect 386848 471454 387168 471486
rect 386848 471218 386890 471454
rect 387126 471218 387168 471454
rect 386848 471134 387168 471218
rect 386848 470898 386890 471134
rect 387126 470898 387168 471134
rect 386848 470866 387168 470898
rect 417568 471454 417888 471486
rect 417568 471218 417610 471454
rect 417846 471218 417888 471454
rect 417568 471134 417888 471218
rect 417568 470898 417610 471134
rect 417846 470898 417888 471134
rect 417568 470866 417888 470898
rect 448288 471454 448608 471486
rect 448288 471218 448330 471454
rect 448566 471218 448608 471454
rect 448288 471134 448608 471218
rect 448288 470898 448330 471134
rect 448566 470898 448608 471134
rect 448288 470866 448608 470898
rect 479008 471454 479328 471486
rect 479008 471218 479050 471454
rect 479286 471218 479328 471454
rect 479008 471134 479328 471218
rect 479008 470898 479050 471134
rect 479286 470898 479328 471134
rect 479008 470866 479328 470898
rect 509728 471454 510048 471486
rect 509728 471218 509770 471454
rect 510006 471218 510048 471454
rect 509728 471134 510048 471218
rect 509728 470898 509770 471134
rect 510006 470898 510048 471134
rect 509728 470866 510048 470898
rect 540448 471454 540768 471486
rect 540448 471218 540490 471454
rect 540726 471218 540768 471454
rect 540448 471134 540768 471218
rect 540448 470898 540490 471134
rect 540726 470898 540768 471134
rect 540448 470866 540768 470898
rect 33568 453454 33888 453486
rect 33568 453218 33610 453454
rect 33846 453218 33888 453454
rect 33568 453134 33888 453218
rect 33568 452898 33610 453134
rect 33846 452898 33888 453134
rect 33568 452866 33888 452898
rect 64288 453454 64608 453486
rect 64288 453218 64330 453454
rect 64566 453218 64608 453454
rect 64288 453134 64608 453218
rect 64288 452898 64330 453134
rect 64566 452898 64608 453134
rect 64288 452866 64608 452898
rect 95008 453454 95328 453486
rect 95008 453218 95050 453454
rect 95286 453218 95328 453454
rect 95008 453134 95328 453218
rect 95008 452898 95050 453134
rect 95286 452898 95328 453134
rect 95008 452866 95328 452898
rect 125728 453454 126048 453486
rect 125728 453218 125770 453454
rect 126006 453218 126048 453454
rect 125728 453134 126048 453218
rect 125728 452898 125770 453134
rect 126006 452898 126048 453134
rect 125728 452866 126048 452898
rect 156448 453454 156768 453486
rect 156448 453218 156490 453454
rect 156726 453218 156768 453454
rect 156448 453134 156768 453218
rect 156448 452898 156490 453134
rect 156726 452898 156768 453134
rect 156448 452866 156768 452898
rect 187168 453454 187488 453486
rect 187168 453218 187210 453454
rect 187446 453218 187488 453454
rect 187168 453134 187488 453218
rect 187168 452898 187210 453134
rect 187446 452898 187488 453134
rect 187168 452866 187488 452898
rect 217888 453454 218208 453486
rect 217888 453218 217930 453454
rect 218166 453218 218208 453454
rect 217888 453134 218208 453218
rect 217888 452898 217930 453134
rect 218166 452898 218208 453134
rect 217888 452866 218208 452898
rect 248608 453454 248928 453486
rect 248608 453218 248650 453454
rect 248886 453218 248928 453454
rect 248608 453134 248928 453218
rect 248608 452898 248650 453134
rect 248886 452898 248928 453134
rect 248608 452866 248928 452898
rect 279328 453454 279648 453486
rect 279328 453218 279370 453454
rect 279606 453218 279648 453454
rect 279328 453134 279648 453218
rect 279328 452898 279370 453134
rect 279606 452898 279648 453134
rect 279328 452866 279648 452898
rect 310048 453454 310368 453486
rect 310048 453218 310090 453454
rect 310326 453218 310368 453454
rect 310048 453134 310368 453218
rect 310048 452898 310090 453134
rect 310326 452898 310368 453134
rect 310048 452866 310368 452898
rect 340768 453454 341088 453486
rect 340768 453218 340810 453454
rect 341046 453218 341088 453454
rect 340768 453134 341088 453218
rect 340768 452898 340810 453134
rect 341046 452898 341088 453134
rect 340768 452866 341088 452898
rect 371488 453454 371808 453486
rect 371488 453218 371530 453454
rect 371766 453218 371808 453454
rect 371488 453134 371808 453218
rect 371488 452898 371530 453134
rect 371766 452898 371808 453134
rect 371488 452866 371808 452898
rect 402208 453454 402528 453486
rect 402208 453218 402250 453454
rect 402486 453218 402528 453454
rect 402208 453134 402528 453218
rect 402208 452898 402250 453134
rect 402486 452898 402528 453134
rect 402208 452866 402528 452898
rect 432928 453454 433248 453486
rect 432928 453218 432970 453454
rect 433206 453218 433248 453454
rect 432928 453134 433248 453218
rect 432928 452898 432970 453134
rect 433206 452898 433248 453134
rect 432928 452866 433248 452898
rect 463648 453454 463968 453486
rect 463648 453218 463690 453454
rect 463926 453218 463968 453454
rect 463648 453134 463968 453218
rect 463648 452898 463690 453134
rect 463926 452898 463968 453134
rect 463648 452866 463968 452898
rect 494368 453454 494688 453486
rect 494368 453218 494410 453454
rect 494646 453218 494688 453454
rect 494368 453134 494688 453218
rect 494368 452898 494410 453134
rect 494646 452898 494688 453134
rect 494368 452866 494688 452898
rect 525088 453454 525408 453486
rect 525088 453218 525130 453454
rect 525366 453218 525408 453454
rect 525088 453134 525408 453218
rect 525088 452898 525130 453134
rect 525366 452898 525408 453134
rect 525088 452866 525408 452898
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 18208 435454 18528 435486
rect 18208 435218 18250 435454
rect 18486 435218 18528 435454
rect 18208 435134 18528 435218
rect 18208 434898 18250 435134
rect 18486 434898 18528 435134
rect 18208 434866 18528 434898
rect 48928 435454 49248 435486
rect 48928 435218 48970 435454
rect 49206 435218 49248 435454
rect 48928 435134 49248 435218
rect 48928 434898 48970 435134
rect 49206 434898 49248 435134
rect 48928 434866 49248 434898
rect 79648 435454 79968 435486
rect 79648 435218 79690 435454
rect 79926 435218 79968 435454
rect 79648 435134 79968 435218
rect 79648 434898 79690 435134
rect 79926 434898 79968 435134
rect 79648 434866 79968 434898
rect 110368 435454 110688 435486
rect 110368 435218 110410 435454
rect 110646 435218 110688 435454
rect 110368 435134 110688 435218
rect 110368 434898 110410 435134
rect 110646 434898 110688 435134
rect 110368 434866 110688 434898
rect 141088 435454 141408 435486
rect 141088 435218 141130 435454
rect 141366 435218 141408 435454
rect 141088 435134 141408 435218
rect 141088 434898 141130 435134
rect 141366 434898 141408 435134
rect 141088 434866 141408 434898
rect 171808 435454 172128 435486
rect 171808 435218 171850 435454
rect 172086 435218 172128 435454
rect 171808 435134 172128 435218
rect 171808 434898 171850 435134
rect 172086 434898 172128 435134
rect 171808 434866 172128 434898
rect 202528 435454 202848 435486
rect 202528 435218 202570 435454
rect 202806 435218 202848 435454
rect 202528 435134 202848 435218
rect 202528 434898 202570 435134
rect 202806 434898 202848 435134
rect 202528 434866 202848 434898
rect 233248 435454 233568 435486
rect 233248 435218 233290 435454
rect 233526 435218 233568 435454
rect 233248 435134 233568 435218
rect 233248 434898 233290 435134
rect 233526 434898 233568 435134
rect 233248 434866 233568 434898
rect 263968 435454 264288 435486
rect 263968 435218 264010 435454
rect 264246 435218 264288 435454
rect 263968 435134 264288 435218
rect 263968 434898 264010 435134
rect 264246 434898 264288 435134
rect 263968 434866 264288 434898
rect 294688 435454 295008 435486
rect 294688 435218 294730 435454
rect 294966 435218 295008 435454
rect 294688 435134 295008 435218
rect 294688 434898 294730 435134
rect 294966 434898 295008 435134
rect 294688 434866 295008 434898
rect 325408 435454 325728 435486
rect 325408 435218 325450 435454
rect 325686 435218 325728 435454
rect 325408 435134 325728 435218
rect 325408 434898 325450 435134
rect 325686 434898 325728 435134
rect 325408 434866 325728 434898
rect 356128 435454 356448 435486
rect 356128 435218 356170 435454
rect 356406 435218 356448 435454
rect 356128 435134 356448 435218
rect 356128 434898 356170 435134
rect 356406 434898 356448 435134
rect 356128 434866 356448 434898
rect 386848 435454 387168 435486
rect 386848 435218 386890 435454
rect 387126 435218 387168 435454
rect 386848 435134 387168 435218
rect 386848 434898 386890 435134
rect 387126 434898 387168 435134
rect 386848 434866 387168 434898
rect 417568 435454 417888 435486
rect 417568 435218 417610 435454
rect 417846 435218 417888 435454
rect 417568 435134 417888 435218
rect 417568 434898 417610 435134
rect 417846 434898 417888 435134
rect 417568 434866 417888 434898
rect 448288 435454 448608 435486
rect 448288 435218 448330 435454
rect 448566 435218 448608 435454
rect 448288 435134 448608 435218
rect 448288 434898 448330 435134
rect 448566 434898 448608 435134
rect 448288 434866 448608 434898
rect 479008 435454 479328 435486
rect 479008 435218 479050 435454
rect 479286 435218 479328 435454
rect 479008 435134 479328 435218
rect 479008 434898 479050 435134
rect 479286 434898 479328 435134
rect 479008 434866 479328 434898
rect 509728 435454 510048 435486
rect 509728 435218 509770 435454
rect 510006 435218 510048 435454
rect 509728 435134 510048 435218
rect 509728 434898 509770 435134
rect 510006 434898 510048 435134
rect 509728 434866 510048 434898
rect 540448 435454 540768 435486
rect 540448 435218 540490 435454
rect 540726 435218 540768 435454
rect 540448 435134 540768 435218
rect 540448 434898 540490 435134
rect 540726 434898 540768 435134
rect 540448 434866 540768 434898
rect 33568 417454 33888 417486
rect 33568 417218 33610 417454
rect 33846 417218 33888 417454
rect 33568 417134 33888 417218
rect 33568 416898 33610 417134
rect 33846 416898 33888 417134
rect 33568 416866 33888 416898
rect 64288 417454 64608 417486
rect 64288 417218 64330 417454
rect 64566 417218 64608 417454
rect 64288 417134 64608 417218
rect 64288 416898 64330 417134
rect 64566 416898 64608 417134
rect 64288 416866 64608 416898
rect 95008 417454 95328 417486
rect 95008 417218 95050 417454
rect 95286 417218 95328 417454
rect 95008 417134 95328 417218
rect 95008 416898 95050 417134
rect 95286 416898 95328 417134
rect 95008 416866 95328 416898
rect 125728 417454 126048 417486
rect 125728 417218 125770 417454
rect 126006 417218 126048 417454
rect 125728 417134 126048 417218
rect 125728 416898 125770 417134
rect 126006 416898 126048 417134
rect 125728 416866 126048 416898
rect 156448 417454 156768 417486
rect 156448 417218 156490 417454
rect 156726 417218 156768 417454
rect 156448 417134 156768 417218
rect 156448 416898 156490 417134
rect 156726 416898 156768 417134
rect 156448 416866 156768 416898
rect 187168 417454 187488 417486
rect 187168 417218 187210 417454
rect 187446 417218 187488 417454
rect 187168 417134 187488 417218
rect 187168 416898 187210 417134
rect 187446 416898 187488 417134
rect 187168 416866 187488 416898
rect 217888 417454 218208 417486
rect 217888 417218 217930 417454
rect 218166 417218 218208 417454
rect 217888 417134 218208 417218
rect 217888 416898 217930 417134
rect 218166 416898 218208 417134
rect 217888 416866 218208 416898
rect 248608 417454 248928 417486
rect 248608 417218 248650 417454
rect 248886 417218 248928 417454
rect 248608 417134 248928 417218
rect 248608 416898 248650 417134
rect 248886 416898 248928 417134
rect 248608 416866 248928 416898
rect 279328 417454 279648 417486
rect 279328 417218 279370 417454
rect 279606 417218 279648 417454
rect 279328 417134 279648 417218
rect 279328 416898 279370 417134
rect 279606 416898 279648 417134
rect 279328 416866 279648 416898
rect 310048 417454 310368 417486
rect 310048 417218 310090 417454
rect 310326 417218 310368 417454
rect 310048 417134 310368 417218
rect 310048 416898 310090 417134
rect 310326 416898 310368 417134
rect 310048 416866 310368 416898
rect 340768 417454 341088 417486
rect 340768 417218 340810 417454
rect 341046 417218 341088 417454
rect 340768 417134 341088 417218
rect 340768 416898 340810 417134
rect 341046 416898 341088 417134
rect 340768 416866 341088 416898
rect 371488 417454 371808 417486
rect 371488 417218 371530 417454
rect 371766 417218 371808 417454
rect 371488 417134 371808 417218
rect 371488 416898 371530 417134
rect 371766 416898 371808 417134
rect 371488 416866 371808 416898
rect 402208 417454 402528 417486
rect 402208 417218 402250 417454
rect 402486 417218 402528 417454
rect 402208 417134 402528 417218
rect 402208 416898 402250 417134
rect 402486 416898 402528 417134
rect 402208 416866 402528 416898
rect 432928 417454 433248 417486
rect 432928 417218 432970 417454
rect 433206 417218 433248 417454
rect 432928 417134 433248 417218
rect 432928 416898 432970 417134
rect 433206 416898 433248 417134
rect 432928 416866 433248 416898
rect 463648 417454 463968 417486
rect 463648 417218 463690 417454
rect 463926 417218 463968 417454
rect 463648 417134 463968 417218
rect 463648 416898 463690 417134
rect 463926 416898 463968 417134
rect 463648 416866 463968 416898
rect 494368 417454 494688 417486
rect 494368 417218 494410 417454
rect 494646 417218 494688 417454
rect 494368 417134 494688 417218
rect 494368 416898 494410 417134
rect 494646 416898 494688 417134
rect 494368 416866 494688 416898
rect 525088 417454 525408 417486
rect 525088 417218 525130 417454
rect 525366 417218 525408 417454
rect 525088 417134 525408 417218
rect 525088 416898 525130 417134
rect 525366 416898 525408 417134
rect 525088 416866 525408 416898
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 18208 399454 18528 399486
rect 18208 399218 18250 399454
rect 18486 399218 18528 399454
rect 18208 399134 18528 399218
rect 18208 398898 18250 399134
rect 18486 398898 18528 399134
rect 18208 398866 18528 398898
rect 48928 399454 49248 399486
rect 48928 399218 48970 399454
rect 49206 399218 49248 399454
rect 48928 399134 49248 399218
rect 48928 398898 48970 399134
rect 49206 398898 49248 399134
rect 48928 398866 49248 398898
rect 79648 399454 79968 399486
rect 79648 399218 79690 399454
rect 79926 399218 79968 399454
rect 79648 399134 79968 399218
rect 79648 398898 79690 399134
rect 79926 398898 79968 399134
rect 79648 398866 79968 398898
rect 110368 399454 110688 399486
rect 110368 399218 110410 399454
rect 110646 399218 110688 399454
rect 110368 399134 110688 399218
rect 110368 398898 110410 399134
rect 110646 398898 110688 399134
rect 110368 398866 110688 398898
rect 141088 399454 141408 399486
rect 141088 399218 141130 399454
rect 141366 399218 141408 399454
rect 141088 399134 141408 399218
rect 141088 398898 141130 399134
rect 141366 398898 141408 399134
rect 141088 398866 141408 398898
rect 171808 399454 172128 399486
rect 171808 399218 171850 399454
rect 172086 399218 172128 399454
rect 171808 399134 172128 399218
rect 171808 398898 171850 399134
rect 172086 398898 172128 399134
rect 171808 398866 172128 398898
rect 202528 399454 202848 399486
rect 202528 399218 202570 399454
rect 202806 399218 202848 399454
rect 202528 399134 202848 399218
rect 202528 398898 202570 399134
rect 202806 398898 202848 399134
rect 202528 398866 202848 398898
rect 233248 399454 233568 399486
rect 233248 399218 233290 399454
rect 233526 399218 233568 399454
rect 233248 399134 233568 399218
rect 233248 398898 233290 399134
rect 233526 398898 233568 399134
rect 233248 398866 233568 398898
rect 263968 399454 264288 399486
rect 263968 399218 264010 399454
rect 264246 399218 264288 399454
rect 263968 399134 264288 399218
rect 263968 398898 264010 399134
rect 264246 398898 264288 399134
rect 263968 398866 264288 398898
rect 294688 399454 295008 399486
rect 294688 399218 294730 399454
rect 294966 399218 295008 399454
rect 294688 399134 295008 399218
rect 294688 398898 294730 399134
rect 294966 398898 295008 399134
rect 294688 398866 295008 398898
rect 325408 399454 325728 399486
rect 325408 399218 325450 399454
rect 325686 399218 325728 399454
rect 325408 399134 325728 399218
rect 325408 398898 325450 399134
rect 325686 398898 325728 399134
rect 325408 398866 325728 398898
rect 356128 399454 356448 399486
rect 356128 399218 356170 399454
rect 356406 399218 356448 399454
rect 356128 399134 356448 399218
rect 356128 398898 356170 399134
rect 356406 398898 356448 399134
rect 356128 398866 356448 398898
rect 386848 399454 387168 399486
rect 386848 399218 386890 399454
rect 387126 399218 387168 399454
rect 386848 399134 387168 399218
rect 386848 398898 386890 399134
rect 387126 398898 387168 399134
rect 386848 398866 387168 398898
rect 417568 399454 417888 399486
rect 417568 399218 417610 399454
rect 417846 399218 417888 399454
rect 417568 399134 417888 399218
rect 417568 398898 417610 399134
rect 417846 398898 417888 399134
rect 417568 398866 417888 398898
rect 448288 399454 448608 399486
rect 448288 399218 448330 399454
rect 448566 399218 448608 399454
rect 448288 399134 448608 399218
rect 448288 398898 448330 399134
rect 448566 398898 448608 399134
rect 448288 398866 448608 398898
rect 479008 399454 479328 399486
rect 479008 399218 479050 399454
rect 479286 399218 479328 399454
rect 479008 399134 479328 399218
rect 479008 398898 479050 399134
rect 479286 398898 479328 399134
rect 479008 398866 479328 398898
rect 509728 399454 510048 399486
rect 509728 399218 509770 399454
rect 510006 399218 510048 399454
rect 509728 399134 510048 399218
rect 509728 398898 509770 399134
rect 510006 398898 510048 399134
rect 509728 398866 510048 398898
rect 540448 399454 540768 399486
rect 540448 399218 540490 399454
rect 540726 399218 540768 399454
rect 540448 399134 540768 399218
rect 540448 398898 540490 399134
rect 540726 398898 540768 399134
rect 540448 398866 540768 398898
rect 33568 381454 33888 381486
rect 33568 381218 33610 381454
rect 33846 381218 33888 381454
rect 33568 381134 33888 381218
rect 33568 380898 33610 381134
rect 33846 380898 33888 381134
rect 33568 380866 33888 380898
rect 64288 381454 64608 381486
rect 64288 381218 64330 381454
rect 64566 381218 64608 381454
rect 64288 381134 64608 381218
rect 64288 380898 64330 381134
rect 64566 380898 64608 381134
rect 64288 380866 64608 380898
rect 95008 381454 95328 381486
rect 95008 381218 95050 381454
rect 95286 381218 95328 381454
rect 95008 381134 95328 381218
rect 95008 380898 95050 381134
rect 95286 380898 95328 381134
rect 95008 380866 95328 380898
rect 125728 381454 126048 381486
rect 125728 381218 125770 381454
rect 126006 381218 126048 381454
rect 125728 381134 126048 381218
rect 125728 380898 125770 381134
rect 126006 380898 126048 381134
rect 125728 380866 126048 380898
rect 156448 381454 156768 381486
rect 156448 381218 156490 381454
rect 156726 381218 156768 381454
rect 156448 381134 156768 381218
rect 156448 380898 156490 381134
rect 156726 380898 156768 381134
rect 156448 380866 156768 380898
rect 187168 381454 187488 381486
rect 187168 381218 187210 381454
rect 187446 381218 187488 381454
rect 187168 381134 187488 381218
rect 187168 380898 187210 381134
rect 187446 380898 187488 381134
rect 187168 380866 187488 380898
rect 217888 381454 218208 381486
rect 217888 381218 217930 381454
rect 218166 381218 218208 381454
rect 217888 381134 218208 381218
rect 217888 380898 217930 381134
rect 218166 380898 218208 381134
rect 217888 380866 218208 380898
rect 248608 381454 248928 381486
rect 248608 381218 248650 381454
rect 248886 381218 248928 381454
rect 248608 381134 248928 381218
rect 248608 380898 248650 381134
rect 248886 380898 248928 381134
rect 248608 380866 248928 380898
rect 279328 381454 279648 381486
rect 279328 381218 279370 381454
rect 279606 381218 279648 381454
rect 279328 381134 279648 381218
rect 279328 380898 279370 381134
rect 279606 380898 279648 381134
rect 279328 380866 279648 380898
rect 310048 381454 310368 381486
rect 310048 381218 310090 381454
rect 310326 381218 310368 381454
rect 310048 381134 310368 381218
rect 310048 380898 310090 381134
rect 310326 380898 310368 381134
rect 310048 380866 310368 380898
rect 340768 381454 341088 381486
rect 340768 381218 340810 381454
rect 341046 381218 341088 381454
rect 340768 381134 341088 381218
rect 340768 380898 340810 381134
rect 341046 380898 341088 381134
rect 340768 380866 341088 380898
rect 371488 381454 371808 381486
rect 371488 381218 371530 381454
rect 371766 381218 371808 381454
rect 371488 381134 371808 381218
rect 371488 380898 371530 381134
rect 371766 380898 371808 381134
rect 371488 380866 371808 380898
rect 402208 381454 402528 381486
rect 402208 381218 402250 381454
rect 402486 381218 402528 381454
rect 402208 381134 402528 381218
rect 402208 380898 402250 381134
rect 402486 380898 402528 381134
rect 402208 380866 402528 380898
rect 432928 381454 433248 381486
rect 432928 381218 432970 381454
rect 433206 381218 433248 381454
rect 432928 381134 433248 381218
rect 432928 380898 432970 381134
rect 433206 380898 433248 381134
rect 432928 380866 433248 380898
rect 463648 381454 463968 381486
rect 463648 381218 463690 381454
rect 463926 381218 463968 381454
rect 463648 381134 463968 381218
rect 463648 380898 463690 381134
rect 463926 380898 463968 381134
rect 463648 380866 463968 380898
rect 494368 381454 494688 381486
rect 494368 381218 494410 381454
rect 494646 381218 494688 381454
rect 494368 381134 494688 381218
rect 494368 380898 494410 381134
rect 494646 380898 494688 381134
rect 494368 380866 494688 380898
rect 525088 381454 525408 381486
rect 525088 381218 525130 381454
rect 525366 381218 525408 381454
rect 525088 381134 525408 381218
rect 525088 380898 525130 381134
rect 525366 380898 525408 381134
rect 525088 380866 525408 380898
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 18208 363454 18528 363486
rect 18208 363218 18250 363454
rect 18486 363218 18528 363454
rect 18208 363134 18528 363218
rect 18208 362898 18250 363134
rect 18486 362898 18528 363134
rect 18208 362866 18528 362898
rect 48928 363454 49248 363486
rect 48928 363218 48970 363454
rect 49206 363218 49248 363454
rect 48928 363134 49248 363218
rect 48928 362898 48970 363134
rect 49206 362898 49248 363134
rect 48928 362866 49248 362898
rect 79648 363454 79968 363486
rect 79648 363218 79690 363454
rect 79926 363218 79968 363454
rect 79648 363134 79968 363218
rect 79648 362898 79690 363134
rect 79926 362898 79968 363134
rect 79648 362866 79968 362898
rect 110368 363454 110688 363486
rect 110368 363218 110410 363454
rect 110646 363218 110688 363454
rect 110368 363134 110688 363218
rect 110368 362898 110410 363134
rect 110646 362898 110688 363134
rect 110368 362866 110688 362898
rect 141088 363454 141408 363486
rect 141088 363218 141130 363454
rect 141366 363218 141408 363454
rect 141088 363134 141408 363218
rect 141088 362898 141130 363134
rect 141366 362898 141408 363134
rect 141088 362866 141408 362898
rect 171808 363454 172128 363486
rect 171808 363218 171850 363454
rect 172086 363218 172128 363454
rect 171808 363134 172128 363218
rect 171808 362898 171850 363134
rect 172086 362898 172128 363134
rect 171808 362866 172128 362898
rect 202528 363454 202848 363486
rect 202528 363218 202570 363454
rect 202806 363218 202848 363454
rect 202528 363134 202848 363218
rect 202528 362898 202570 363134
rect 202806 362898 202848 363134
rect 202528 362866 202848 362898
rect 233248 363454 233568 363486
rect 233248 363218 233290 363454
rect 233526 363218 233568 363454
rect 233248 363134 233568 363218
rect 233248 362898 233290 363134
rect 233526 362898 233568 363134
rect 233248 362866 233568 362898
rect 263968 363454 264288 363486
rect 263968 363218 264010 363454
rect 264246 363218 264288 363454
rect 263968 363134 264288 363218
rect 263968 362898 264010 363134
rect 264246 362898 264288 363134
rect 263968 362866 264288 362898
rect 294688 363454 295008 363486
rect 294688 363218 294730 363454
rect 294966 363218 295008 363454
rect 294688 363134 295008 363218
rect 294688 362898 294730 363134
rect 294966 362898 295008 363134
rect 294688 362866 295008 362898
rect 325408 363454 325728 363486
rect 325408 363218 325450 363454
rect 325686 363218 325728 363454
rect 325408 363134 325728 363218
rect 325408 362898 325450 363134
rect 325686 362898 325728 363134
rect 325408 362866 325728 362898
rect 356128 363454 356448 363486
rect 356128 363218 356170 363454
rect 356406 363218 356448 363454
rect 356128 363134 356448 363218
rect 356128 362898 356170 363134
rect 356406 362898 356448 363134
rect 356128 362866 356448 362898
rect 386848 363454 387168 363486
rect 386848 363218 386890 363454
rect 387126 363218 387168 363454
rect 386848 363134 387168 363218
rect 386848 362898 386890 363134
rect 387126 362898 387168 363134
rect 386848 362866 387168 362898
rect 417568 363454 417888 363486
rect 417568 363218 417610 363454
rect 417846 363218 417888 363454
rect 417568 363134 417888 363218
rect 417568 362898 417610 363134
rect 417846 362898 417888 363134
rect 417568 362866 417888 362898
rect 448288 363454 448608 363486
rect 448288 363218 448330 363454
rect 448566 363218 448608 363454
rect 448288 363134 448608 363218
rect 448288 362898 448330 363134
rect 448566 362898 448608 363134
rect 448288 362866 448608 362898
rect 479008 363454 479328 363486
rect 479008 363218 479050 363454
rect 479286 363218 479328 363454
rect 479008 363134 479328 363218
rect 479008 362898 479050 363134
rect 479286 362898 479328 363134
rect 479008 362866 479328 362898
rect 509728 363454 510048 363486
rect 509728 363218 509770 363454
rect 510006 363218 510048 363454
rect 509728 363134 510048 363218
rect 509728 362898 509770 363134
rect 510006 362898 510048 363134
rect 509728 362866 510048 362898
rect 540448 363454 540768 363486
rect 540448 363218 540490 363454
rect 540726 363218 540768 363454
rect 540448 363134 540768 363218
rect 540448 362898 540490 363134
rect 540726 362898 540768 363134
rect 540448 362866 540768 362898
rect 33568 345454 33888 345486
rect 33568 345218 33610 345454
rect 33846 345218 33888 345454
rect 33568 345134 33888 345218
rect 33568 344898 33610 345134
rect 33846 344898 33888 345134
rect 33568 344866 33888 344898
rect 64288 345454 64608 345486
rect 64288 345218 64330 345454
rect 64566 345218 64608 345454
rect 64288 345134 64608 345218
rect 64288 344898 64330 345134
rect 64566 344898 64608 345134
rect 64288 344866 64608 344898
rect 95008 345454 95328 345486
rect 95008 345218 95050 345454
rect 95286 345218 95328 345454
rect 95008 345134 95328 345218
rect 95008 344898 95050 345134
rect 95286 344898 95328 345134
rect 95008 344866 95328 344898
rect 125728 345454 126048 345486
rect 125728 345218 125770 345454
rect 126006 345218 126048 345454
rect 125728 345134 126048 345218
rect 125728 344898 125770 345134
rect 126006 344898 126048 345134
rect 125728 344866 126048 344898
rect 156448 345454 156768 345486
rect 156448 345218 156490 345454
rect 156726 345218 156768 345454
rect 156448 345134 156768 345218
rect 156448 344898 156490 345134
rect 156726 344898 156768 345134
rect 156448 344866 156768 344898
rect 187168 345454 187488 345486
rect 187168 345218 187210 345454
rect 187446 345218 187488 345454
rect 187168 345134 187488 345218
rect 187168 344898 187210 345134
rect 187446 344898 187488 345134
rect 187168 344866 187488 344898
rect 217888 345454 218208 345486
rect 217888 345218 217930 345454
rect 218166 345218 218208 345454
rect 217888 345134 218208 345218
rect 217888 344898 217930 345134
rect 218166 344898 218208 345134
rect 217888 344866 218208 344898
rect 248608 345454 248928 345486
rect 248608 345218 248650 345454
rect 248886 345218 248928 345454
rect 248608 345134 248928 345218
rect 248608 344898 248650 345134
rect 248886 344898 248928 345134
rect 248608 344866 248928 344898
rect 279328 345454 279648 345486
rect 279328 345218 279370 345454
rect 279606 345218 279648 345454
rect 279328 345134 279648 345218
rect 279328 344898 279370 345134
rect 279606 344898 279648 345134
rect 279328 344866 279648 344898
rect 310048 345454 310368 345486
rect 310048 345218 310090 345454
rect 310326 345218 310368 345454
rect 310048 345134 310368 345218
rect 310048 344898 310090 345134
rect 310326 344898 310368 345134
rect 310048 344866 310368 344898
rect 340768 345454 341088 345486
rect 340768 345218 340810 345454
rect 341046 345218 341088 345454
rect 340768 345134 341088 345218
rect 340768 344898 340810 345134
rect 341046 344898 341088 345134
rect 340768 344866 341088 344898
rect 371488 345454 371808 345486
rect 371488 345218 371530 345454
rect 371766 345218 371808 345454
rect 371488 345134 371808 345218
rect 371488 344898 371530 345134
rect 371766 344898 371808 345134
rect 371488 344866 371808 344898
rect 402208 345454 402528 345486
rect 402208 345218 402250 345454
rect 402486 345218 402528 345454
rect 402208 345134 402528 345218
rect 402208 344898 402250 345134
rect 402486 344898 402528 345134
rect 402208 344866 402528 344898
rect 432928 345454 433248 345486
rect 432928 345218 432970 345454
rect 433206 345218 433248 345454
rect 432928 345134 433248 345218
rect 432928 344898 432970 345134
rect 433206 344898 433248 345134
rect 432928 344866 433248 344898
rect 463648 345454 463968 345486
rect 463648 345218 463690 345454
rect 463926 345218 463968 345454
rect 463648 345134 463968 345218
rect 463648 344898 463690 345134
rect 463926 344898 463968 345134
rect 463648 344866 463968 344898
rect 494368 345454 494688 345486
rect 494368 345218 494410 345454
rect 494646 345218 494688 345454
rect 494368 345134 494688 345218
rect 494368 344898 494410 345134
rect 494646 344898 494688 345134
rect 494368 344866 494688 344898
rect 525088 345454 525408 345486
rect 525088 345218 525130 345454
rect 525366 345218 525408 345454
rect 525088 345134 525408 345218
rect 525088 344898 525130 345134
rect 525366 344898 525408 345134
rect 525088 344866 525408 344898
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 18208 327454 18528 327486
rect 18208 327218 18250 327454
rect 18486 327218 18528 327454
rect 18208 327134 18528 327218
rect 18208 326898 18250 327134
rect 18486 326898 18528 327134
rect 18208 326866 18528 326898
rect 48928 327454 49248 327486
rect 48928 327218 48970 327454
rect 49206 327218 49248 327454
rect 48928 327134 49248 327218
rect 48928 326898 48970 327134
rect 49206 326898 49248 327134
rect 48928 326866 49248 326898
rect 79648 327454 79968 327486
rect 79648 327218 79690 327454
rect 79926 327218 79968 327454
rect 79648 327134 79968 327218
rect 79648 326898 79690 327134
rect 79926 326898 79968 327134
rect 79648 326866 79968 326898
rect 110368 327454 110688 327486
rect 110368 327218 110410 327454
rect 110646 327218 110688 327454
rect 110368 327134 110688 327218
rect 110368 326898 110410 327134
rect 110646 326898 110688 327134
rect 110368 326866 110688 326898
rect 141088 327454 141408 327486
rect 141088 327218 141130 327454
rect 141366 327218 141408 327454
rect 141088 327134 141408 327218
rect 141088 326898 141130 327134
rect 141366 326898 141408 327134
rect 141088 326866 141408 326898
rect 171808 327454 172128 327486
rect 171808 327218 171850 327454
rect 172086 327218 172128 327454
rect 171808 327134 172128 327218
rect 171808 326898 171850 327134
rect 172086 326898 172128 327134
rect 171808 326866 172128 326898
rect 202528 327454 202848 327486
rect 202528 327218 202570 327454
rect 202806 327218 202848 327454
rect 202528 327134 202848 327218
rect 202528 326898 202570 327134
rect 202806 326898 202848 327134
rect 202528 326866 202848 326898
rect 233248 327454 233568 327486
rect 233248 327218 233290 327454
rect 233526 327218 233568 327454
rect 233248 327134 233568 327218
rect 233248 326898 233290 327134
rect 233526 326898 233568 327134
rect 233248 326866 233568 326898
rect 263968 327454 264288 327486
rect 263968 327218 264010 327454
rect 264246 327218 264288 327454
rect 263968 327134 264288 327218
rect 263968 326898 264010 327134
rect 264246 326898 264288 327134
rect 263968 326866 264288 326898
rect 294688 327454 295008 327486
rect 294688 327218 294730 327454
rect 294966 327218 295008 327454
rect 294688 327134 295008 327218
rect 294688 326898 294730 327134
rect 294966 326898 295008 327134
rect 294688 326866 295008 326898
rect 325408 327454 325728 327486
rect 325408 327218 325450 327454
rect 325686 327218 325728 327454
rect 325408 327134 325728 327218
rect 325408 326898 325450 327134
rect 325686 326898 325728 327134
rect 325408 326866 325728 326898
rect 356128 327454 356448 327486
rect 356128 327218 356170 327454
rect 356406 327218 356448 327454
rect 356128 327134 356448 327218
rect 356128 326898 356170 327134
rect 356406 326898 356448 327134
rect 356128 326866 356448 326898
rect 386848 327454 387168 327486
rect 386848 327218 386890 327454
rect 387126 327218 387168 327454
rect 386848 327134 387168 327218
rect 386848 326898 386890 327134
rect 387126 326898 387168 327134
rect 386848 326866 387168 326898
rect 417568 327454 417888 327486
rect 417568 327218 417610 327454
rect 417846 327218 417888 327454
rect 417568 327134 417888 327218
rect 417568 326898 417610 327134
rect 417846 326898 417888 327134
rect 417568 326866 417888 326898
rect 448288 327454 448608 327486
rect 448288 327218 448330 327454
rect 448566 327218 448608 327454
rect 448288 327134 448608 327218
rect 448288 326898 448330 327134
rect 448566 326898 448608 327134
rect 448288 326866 448608 326898
rect 479008 327454 479328 327486
rect 479008 327218 479050 327454
rect 479286 327218 479328 327454
rect 479008 327134 479328 327218
rect 479008 326898 479050 327134
rect 479286 326898 479328 327134
rect 479008 326866 479328 326898
rect 509728 327454 510048 327486
rect 509728 327218 509770 327454
rect 510006 327218 510048 327454
rect 509728 327134 510048 327218
rect 509728 326898 509770 327134
rect 510006 326898 510048 327134
rect 509728 326866 510048 326898
rect 540448 327454 540768 327486
rect 540448 327218 540490 327454
rect 540726 327218 540768 327454
rect 540448 327134 540768 327218
rect 540448 326898 540490 327134
rect 540726 326898 540768 327134
rect 540448 326866 540768 326898
rect 33568 309454 33888 309486
rect 33568 309218 33610 309454
rect 33846 309218 33888 309454
rect 33568 309134 33888 309218
rect 33568 308898 33610 309134
rect 33846 308898 33888 309134
rect 33568 308866 33888 308898
rect 64288 309454 64608 309486
rect 64288 309218 64330 309454
rect 64566 309218 64608 309454
rect 64288 309134 64608 309218
rect 64288 308898 64330 309134
rect 64566 308898 64608 309134
rect 64288 308866 64608 308898
rect 95008 309454 95328 309486
rect 95008 309218 95050 309454
rect 95286 309218 95328 309454
rect 95008 309134 95328 309218
rect 95008 308898 95050 309134
rect 95286 308898 95328 309134
rect 95008 308866 95328 308898
rect 125728 309454 126048 309486
rect 125728 309218 125770 309454
rect 126006 309218 126048 309454
rect 125728 309134 126048 309218
rect 125728 308898 125770 309134
rect 126006 308898 126048 309134
rect 125728 308866 126048 308898
rect 156448 309454 156768 309486
rect 156448 309218 156490 309454
rect 156726 309218 156768 309454
rect 156448 309134 156768 309218
rect 156448 308898 156490 309134
rect 156726 308898 156768 309134
rect 156448 308866 156768 308898
rect 187168 309454 187488 309486
rect 187168 309218 187210 309454
rect 187446 309218 187488 309454
rect 187168 309134 187488 309218
rect 187168 308898 187210 309134
rect 187446 308898 187488 309134
rect 187168 308866 187488 308898
rect 217888 309454 218208 309486
rect 217888 309218 217930 309454
rect 218166 309218 218208 309454
rect 217888 309134 218208 309218
rect 217888 308898 217930 309134
rect 218166 308898 218208 309134
rect 217888 308866 218208 308898
rect 248608 309454 248928 309486
rect 248608 309218 248650 309454
rect 248886 309218 248928 309454
rect 248608 309134 248928 309218
rect 248608 308898 248650 309134
rect 248886 308898 248928 309134
rect 248608 308866 248928 308898
rect 279328 309454 279648 309486
rect 279328 309218 279370 309454
rect 279606 309218 279648 309454
rect 279328 309134 279648 309218
rect 279328 308898 279370 309134
rect 279606 308898 279648 309134
rect 279328 308866 279648 308898
rect 310048 309454 310368 309486
rect 310048 309218 310090 309454
rect 310326 309218 310368 309454
rect 310048 309134 310368 309218
rect 310048 308898 310090 309134
rect 310326 308898 310368 309134
rect 310048 308866 310368 308898
rect 340768 309454 341088 309486
rect 340768 309218 340810 309454
rect 341046 309218 341088 309454
rect 340768 309134 341088 309218
rect 340768 308898 340810 309134
rect 341046 308898 341088 309134
rect 340768 308866 341088 308898
rect 371488 309454 371808 309486
rect 371488 309218 371530 309454
rect 371766 309218 371808 309454
rect 371488 309134 371808 309218
rect 371488 308898 371530 309134
rect 371766 308898 371808 309134
rect 371488 308866 371808 308898
rect 402208 309454 402528 309486
rect 402208 309218 402250 309454
rect 402486 309218 402528 309454
rect 402208 309134 402528 309218
rect 402208 308898 402250 309134
rect 402486 308898 402528 309134
rect 402208 308866 402528 308898
rect 432928 309454 433248 309486
rect 432928 309218 432970 309454
rect 433206 309218 433248 309454
rect 432928 309134 433248 309218
rect 432928 308898 432970 309134
rect 433206 308898 433248 309134
rect 432928 308866 433248 308898
rect 463648 309454 463968 309486
rect 463648 309218 463690 309454
rect 463926 309218 463968 309454
rect 463648 309134 463968 309218
rect 463648 308898 463690 309134
rect 463926 308898 463968 309134
rect 463648 308866 463968 308898
rect 494368 309454 494688 309486
rect 494368 309218 494410 309454
rect 494646 309218 494688 309454
rect 494368 309134 494688 309218
rect 494368 308898 494410 309134
rect 494646 308898 494688 309134
rect 494368 308866 494688 308898
rect 525088 309454 525408 309486
rect 525088 309218 525130 309454
rect 525366 309218 525408 309454
rect 525088 309134 525408 309218
rect 525088 308898 525130 309134
rect 525366 308898 525408 309134
rect 525088 308866 525408 308898
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 18208 291454 18528 291486
rect 18208 291218 18250 291454
rect 18486 291218 18528 291454
rect 18208 291134 18528 291218
rect 18208 290898 18250 291134
rect 18486 290898 18528 291134
rect 18208 290866 18528 290898
rect 48928 291454 49248 291486
rect 48928 291218 48970 291454
rect 49206 291218 49248 291454
rect 48928 291134 49248 291218
rect 48928 290898 48970 291134
rect 49206 290898 49248 291134
rect 48928 290866 49248 290898
rect 79648 291454 79968 291486
rect 79648 291218 79690 291454
rect 79926 291218 79968 291454
rect 79648 291134 79968 291218
rect 79648 290898 79690 291134
rect 79926 290898 79968 291134
rect 79648 290866 79968 290898
rect 110368 291454 110688 291486
rect 110368 291218 110410 291454
rect 110646 291218 110688 291454
rect 110368 291134 110688 291218
rect 110368 290898 110410 291134
rect 110646 290898 110688 291134
rect 110368 290866 110688 290898
rect 141088 291454 141408 291486
rect 141088 291218 141130 291454
rect 141366 291218 141408 291454
rect 141088 291134 141408 291218
rect 141088 290898 141130 291134
rect 141366 290898 141408 291134
rect 141088 290866 141408 290898
rect 171808 291454 172128 291486
rect 171808 291218 171850 291454
rect 172086 291218 172128 291454
rect 171808 291134 172128 291218
rect 171808 290898 171850 291134
rect 172086 290898 172128 291134
rect 171808 290866 172128 290898
rect 202528 291454 202848 291486
rect 202528 291218 202570 291454
rect 202806 291218 202848 291454
rect 202528 291134 202848 291218
rect 202528 290898 202570 291134
rect 202806 290898 202848 291134
rect 202528 290866 202848 290898
rect 233248 291454 233568 291486
rect 233248 291218 233290 291454
rect 233526 291218 233568 291454
rect 233248 291134 233568 291218
rect 233248 290898 233290 291134
rect 233526 290898 233568 291134
rect 233248 290866 233568 290898
rect 263968 291454 264288 291486
rect 263968 291218 264010 291454
rect 264246 291218 264288 291454
rect 263968 291134 264288 291218
rect 263968 290898 264010 291134
rect 264246 290898 264288 291134
rect 263968 290866 264288 290898
rect 294688 291454 295008 291486
rect 294688 291218 294730 291454
rect 294966 291218 295008 291454
rect 294688 291134 295008 291218
rect 294688 290898 294730 291134
rect 294966 290898 295008 291134
rect 294688 290866 295008 290898
rect 325408 291454 325728 291486
rect 325408 291218 325450 291454
rect 325686 291218 325728 291454
rect 325408 291134 325728 291218
rect 325408 290898 325450 291134
rect 325686 290898 325728 291134
rect 325408 290866 325728 290898
rect 356128 291454 356448 291486
rect 356128 291218 356170 291454
rect 356406 291218 356448 291454
rect 356128 291134 356448 291218
rect 356128 290898 356170 291134
rect 356406 290898 356448 291134
rect 356128 290866 356448 290898
rect 386848 291454 387168 291486
rect 386848 291218 386890 291454
rect 387126 291218 387168 291454
rect 386848 291134 387168 291218
rect 386848 290898 386890 291134
rect 387126 290898 387168 291134
rect 386848 290866 387168 290898
rect 417568 291454 417888 291486
rect 417568 291218 417610 291454
rect 417846 291218 417888 291454
rect 417568 291134 417888 291218
rect 417568 290898 417610 291134
rect 417846 290898 417888 291134
rect 417568 290866 417888 290898
rect 448288 291454 448608 291486
rect 448288 291218 448330 291454
rect 448566 291218 448608 291454
rect 448288 291134 448608 291218
rect 448288 290898 448330 291134
rect 448566 290898 448608 291134
rect 448288 290866 448608 290898
rect 479008 291454 479328 291486
rect 479008 291218 479050 291454
rect 479286 291218 479328 291454
rect 479008 291134 479328 291218
rect 479008 290898 479050 291134
rect 479286 290898 479328 291134
rect 479008 290866 479328 290898
rect 509728 291454 510048 291486
rect 509728 291218 509770 291454
rect 510006 291218 510048 291454
rect 509728 291134 510048 291218
rect 509728 290898 509770 291134
rect 510006 290898 510048 291134
rect 509728 290866 510048 290898
rect 540448 291454 540768 291486
rect 540448 291218 540490 291454
rect 540726 291218 540768 291454
rect 540448 291134 540768 291218
rect 540448 290898 540490 291134
rect 540726 290898 540768 291134
rect 540448 290866 540768 290898
rect 33568 273454 33888 273486
rect 33568 273218 33610 273454
rect 33846 273218 33888 273454
rect 33568 273134 33888 273218
rect 33568 272898 33610 273134
rect 33846 272898 33888 273134
rect 33568 272866 33888 272898
rect 64288 273454 64608 273486
rect 64288 273218 64330 273454
rect 64566 273218 64608 273454
rect 64288 273134 64608 273218
rect 64288 272898 64330 273134
rect 64566 272898 64608 273134
rect 64288 272866 64608 272898
rect 95008 273454 95328 273486
rect 95008 273218 95050 273454
rect 95286 273218 95328 273454
rect 95008 273134 95328 273218
rect 95008 272898 95050 273134
rect 95286 272898 95328 273134
rect 95008 272866 95328 272898
rect 125728 273454 126048 273486
rect 125728 273218 125770 273454
rect 126006 273218 126048 273454
rect 125728 273134 126048 273218
rect 125728 272898 125770 273134
rect 126006 272898 126048 273134
rect 125728 272866 126048 272898
rect 156448 273454 156768 273486
rect 156448 273218 156490 273454
rect 156726 273218 156768 273454
rect 156448 273134 156768 273218
rect 156448 272898 156490 273134
rect 156726 272898 156768 273134
rect 156448 272866 156768 272898
rect 187168 273454 187488 273486
rect 187168 273218 187210 273454
rect 187446 273218 187488 273454
rect 187168 273134 187488 273218
rect 187168 272898 187210 273134
rect 187446 272898 187488 273134
rect 187168 272866 187488 272898
rect 217888 273454 218208 273486
rect 217888 273218 217930 273454
rect 218166 273218 218208 273454
rect 217888 273134 218208 273218
rect 217888 272898 217930 273134
rect 218166 272898 218208 273134
rect 217888 272866 218208 272898
rect 248608 273454 248928 273486
rect 248608 273218 248650 273454
rect 248886 273218 248928 273454
rect 248608 273134 248928 273218
rect 248608 272898 248650 273134
rect 248886 272898 248928 273134
rect 248608 272866 248928 272898
rect 279328 273454 279648 273486
rect 279328 273218 279370 273454
rect 279606 273218 279648 273454
rect 279328 273134 279648 273218
rect 279328 272898 279370 273134
rect 279606 272898 279648 273134
rect 279328 272866 279648 272898
rect 310048 273454 310368 273486
rect 310048 273218 310090 273454
rect 310326 273218 310368 273454
rect 310048 273134 310368 273218
rect 310048 272898 310090 273134
rect 310326 272898 310368 273134
rect 310048 272866 310368 272898
rect 340768 273454 341088 273486
rect 340768 273218 340810 273454
rect 341046 273218 341088 273454
rect 340768 273134 341088 273218
rect 340768 272898 340810 273134
rect 341046 272898 341088 273134
rect 340768 272866 341088 272898
rect 371488 273454 371808 273486
rect 371488 273218 371530 273454
rect 371766 273218 371808 273454
rect 371488 273134 371808 273218
rect 371488 272898 371530 273134
rect 371766 272898 371808 273134
rect 371488 272866 371808 272898
rect 402208 273454 402528 273486
rect 402208 273218 402250 273454
rect 402486 273218 402528 273454
rect 402208 273134 402528 273218
rect 402208 272898 402250 273134
rect 402486 272898 402528 273134
rect 402208 272866 402528 272898
rect 432928 273454 433248 273486
rect 432928 273218 432970 273454
rect 433206 273218 433248 273454
rect 432928 273134 433248 273218
rect 432928 272898 432970 273134
rect 433206 272898 433248 273134
rect 432928 272866 433248 272898
rect 463648 273454 463968 273486
rect 463648 273218 463690 273454
rect 463926 273218 463968 273454
rect 463648 273134 463968 273218
rect 463648 272898 463690 273134
rect 463926 272898 463968 273134
rect 463648 272866 463968 272898
rect 494368 273454 494688 273486
rect 494368 273218 494410 273454
rect 494646 273218 494688 273454
rect 494368 273134 494688 273218
rect 494368 272898 494410 273134
rect 494646 272898 494688 273134
rect 494368 272866 494688 272898
rect 525088 273454 525408 273486
rect 525088 273218 525130 273454
rect 525366 273218 525408 273454
rect 525088 273134 525408 273218
rect 525088 272898 525130 273134
rect 525366 272898 525408 273134
rect 525088 272866 525408 272898
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 18208 255454 18528 255486
rect 18208 255218 18250 255454
rect 18486 255218 18528 255454
rect 18208 255134 18528 255218
rect 18208 254898 18250 255134
rect 18486 254898 18528 255134
rect 18208 254866 18528 254898
rect 48928 255454 49248 255486
rect 48928 255218 48970 255454
rect 49206 255218 49248 255454
rect 48928 255134 49248 255218
rect 48928 254898 48970 255134
rect 49206 254898 49248 255134
rect 48928 254866 49248 254898
rect 79648 255454 79968 255486
rect 79648 255218 79690 255454
rect 79926 255218 79968 255454
rect 79648 255134 79968 255218
rect 79648 254898 79690 255134
rect 79926 254898 79968 255134
rect 79648 254866 79968 254898
rect 110368 255454 110688 255486
rect 110368 255218 110410 255454
rect 110646 255218 110688 255454
rect 110368 255134 110688 255218
rect 110368 254898 110410 255134
rect 110646 254898 110688 255134
rect 110368 254866 110688 254898
rect 141088 255454 141408 255486
rect 141088 255218 141130 255454
rect 141366 255218 141408 255454
rect 141088 255134 141408 255218
rect 141088 254898 141130 255134
rect 141366 254898 141408 255134
rect 141088 254866 141408 254898
rect 171808 255454 172128 255486
rect 171808 255218 171850 255454
rect 172086 255218 172128 255454
rect 171808 255134 172128 255218
rect 171808 254898 171850 255134
rect 172086 254898 172128 255134
rect 171808 254866 172128 254898
rect 202528 255454 202848 255486
rect 202528 255218 202570 255454
rect 202806 255218 202848 255454
rect 202528 255134 202848 255218
rect 202528 254898 202570 255134
rect 202806 254898 202848 255134
rect 202528 254866 202848 254898
rect 233248 255454 233568 255486
rect 233248 255218 233290 255454
rect 233526 255218 233568 255454
rect 233248 255134 233568 255218
rect 233248 254898 233290 255134
rect 233526 254898 233568 255134
rect 233248 254866 233568 254898
rect 263968 255454 264288 255486
rect 263968 255218 264010 255454
rect 264246 255218 264288 255454
rect 263968 255134 264288 255218
rect 263968 254898 264010 255134
rect 264246 254898 264288 255134
rect 263968 254866 264288 254898
rect 294688 255454 295008 255486
rect 294688 255218 294730 255454
rect 294966 255218 295008 255454
rect 294688 255134 295008 255218
rect 294688 254898 294730 255134
rect 294966 254898 295008 255134
rect 294688 254866 295008 254898
rect 325408 255454 325728 255486
rect 325408 255218 325450 255454
rect 325686 255218 325728 255454
rect 325408 255134 325728 255218
rect 325408 254898 325450 255134
rect 325686 254898 325728 255134
rect 325408 254866 325728 254898
rect 356128 255454 356448 255486
rect 356128 255218 356170 255454
rect 356406 255218 356448 255454
rect 356128 255134 356448 255218
rect 356128 254898 356170 255134
rect 356406 254898 356448 255134
rect 356128 254866 356448 254898
rect 386848 255454 387168 255486
rect 386848 255218 386890 255454
rect 387126 255218 387168 255454
rect 386848 255134 387168 255218
rect 386848 254898 386890 255134
rect 387126 254898 387168 255134
rect 386848 254866 387168 254898
rect 417568 255454 417888 255486
rect 417568 255218 417610 255454
rect 417846 255218 417888 255454
rect 417568 255134 417888 255218
rect 417568 254898 417610 255134
rect 417846 254898 417888 255134
rect 417568 254866 417888 254898
rect 448288 255454 448608 255486
rect 448288 255218 448330 255454
rect 448566 255218 448608 255454
rect 448288 255134 448608 255218
rect 448288 254898 448330 255134
rect 448566 254898 448608 255134
rect 448288 254866 448608 254898
rect 479008 255454 479328 255486
rect 479008 255218 479050 255454
rect 479286 255218 479328 255454
rect 479008 255134 479328 255218
rect 479008 254898 479050 255134
rect 479286 254898 479328 255134
rect 479008 254866 479328 254898
rect 509728 255454 510048 255486
rect 509728 255218 509770 255454
rect 510006 255218 510048 255454
rect 509728 255134 510048 255218
rect 509728 254898 509770 255134
rect 510006 254898 510048 255134
rect 509728 254866 510048 254898
rect 540448 255454 540768 255486
rect 540448 255218 540490 255454
rect 540726 255218 540768 255454
rect 540448 255134 540768 255218
rect 540448 254898 540490 255134
rect 540726 254898 540768 255134
rect 540448 254866 540768 254898
rect 33568 237454 33888 237486
rect 33568 237218 33610 237454
rect 33846 237218 33888 237454
rect 33568 237134 33888 237218
rect 33568 236898 33610 237134
rect 33846 236898 33888 237134
rect 33568 236866 33888 236898
rect 64288 237454 64608 237486
rect 64288 237218 64330 237454
rect 64566 237218 64608 237454
rect 64288 237134 64608 237218
rect 64288 236898 64330 237134
rect 64566 236898 64608 237134
rect 64288 236866 64608 236898
rect 95008 237454 95328 237486
rect 95008 237218 95050 237454
rect 95286 237218 95328 237454
rect 95008 237134 95328 237218
rect 95008 236898 95050 237134
rect 95286 236898 95328 237134
rect 95008 236866 95328 236898
rect 125728 237454 126048 237486
rect 125728 237218 125770 237454
rect 126006 237218 126048 237454
rect 125728 237134 126048 237218
rect 125728 236898 125770 237134
rect 126006 236898 126048 237134
rect 125728 236866 126048 236898
rect 156448 237454 156768 237486
rect 156448 237218 156490 237454
rect 156726 237218 156768 237454
rect 156448 237134 156768 237218
rect 156448 236898 156490 237134
rect 156726 236898 156768 237134
rect 156448 236866 156768 236898
rect 187168 237454 187488 237486
rect 187168 237218 187210 237454
rect 187446 237218 187488 237454
rect 187168 237134 187488 237218
rect 187168 236898 187210 237134
rect 187446 236898 187488 237134
rect 187168 236866 187488 236898
rect 217888 237454 218208 237486
rect 217888 237218 217930 237454
rect 218166 237218 218208 237454
rect 217888 237134 218208 237218
rect 217888 236898 217930 237134
rect 218166 236898 218208 237134
rect 217888 236866 218208 236898
rect 248608 237454 248928 237486
rect 248608 237218 248650 237454
rect 248886 237218 248928 237454
rect 248608 237134 248928 237218
rect 248608 236898 248650 237134
rect 248886 236898 248928 237134
rect 248608 236866 248928 236898
rect 279328 237454 279648 237486
rect 279328 237218 279370 237454
rect 279606 237218 279648 237454
rect 279328 237134 279648 237218
rect 279328 236898 279370 237134
rect 279606 236898 279648 237134
rect 279328 236866 279648 236898
rect 310048 237454 310368 237486
rect 310048 237218 310090 237454
rect 310326 237218 310368 237454
rect 310048 237134 310368 237218
rect 310048 236898 310090 237134
rect 310326 236898 310368 237134
rect 310048 236866 310368 236898
rect 340768 237454 341088 237486
rect 340768 237218 340810 237454
rect 341046 237218 341088 237454
rect 340768 237134 341088 237218
rect 340768 236898 340810 237134
rect 341046 236898 341088 237134
rect 340768 236866 341088 236898
rect 371488 237454 371808 237486
rect 371488 237218 371530 237454
rect 371766 237218 371808 237454
rect 371488 237134 371808 237218
rect 371488 236898 371530 237134
rect 371766 236898 371808 237134
rect 371488 236866 371808 236898
rect 402208 237454 402528 237486
rect 402208 237218 402250 237454
rect 402486 237218 402528 237454
rect 402208 237134 402528 237218
rect 402208 236898 402250 237134
rect 402486 236898 402528 237134
rect 402208 236866 402528 236898
rect 432928 237454 433248 237486
rect 432928 237218 432970 237454
rect 433206 237218 433248 237454
rect 432928 237134 433248 237218
rect 432928 236898 432970 237134
rect 433206 236898 433248 237134
rect 432928 236866 433248 236898
rect 463648 237454 463968 237486
rect 463648 237218 463690 237454
rect 463926 237218 463968 237454
rect 463648 237134 463968 237218
rect 463648 236898 463690 237134
rect 463926 236898 463968 237134
rect 463648 236866 463968 236898
rect 494368 237454 494688 237486
rect 494368 237218 494410 237454
rect 494646 237218 494688 237454
rect 494368 237134 494688 237218
rect 494368 236898 494410 237134
rect 494646 236898 494688 237134
rect 494368 236866 494688 236898
rect 525088 237454 525408 237486
rect 525088 237218 525130 237454
rect 525366 237218 525408 237454
rect 525088 237134 525408 237218
rect 525088 236898 525130 237134
rect 525366 236898 525408 237134
rect 525088 236866 525408 236898
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 18208 219454 18528 219486
rect 18208 219218 18250 219454
rect 18486 219218 18528 219454
rect 18208 219134 18528 219218
rect 18208 218898 18250 219134
rect 18486 218898 18528 219134
rect 18208 218866 18528 218898
rect 48928 219454 49248 219486
rect 48928 219218 48970 219454
rect 49206 219218 49248 219454
rect 48928 219134 49248 219218
rect 48928 218898 48970 219134
rect 49206 218898 49248 219134
rect 48928 218866 49248 218898
rect 79648 219454 79968 219486
rect 79648 219218 79690 219454
rect 79926 219218 79968 219454
rect 79648 219134 79968 219218
rect 79648 218898 79690 219134
rect 79926 218898 79968 219134
rect 79648 218866 79968 218898
rect 110368 219454 110688 219486
rect 110368 219218 110410 219454
rect 110646 219218 110688 219454
rect 110368 219134 110688 219218
rect 110368 218898 110410 219134
rect 110646 218898 110688 219134
rect 110368 218866 110688 218898
rect 141088 219454 141408 219486
rect 141088 219218 141130 219454
rect 141366 219218 141408 219454
rect 141088 219134 141408 219218
rect 141088 218898 141130 219134
rect 141366 218898 141408 219134
rect 141088 218866 141408 218898
rect 171808 219454 172128 219486
rect 171808 219218 171850 219454
rect 172086 219218 172128 219454
rect 171808 219134 172128 219218
rect 171808 218898 171850 219134
rect 172086 218898 172128 219134
rect 171808 218866 172128 218898
rect 202528 219454 202848 219486
rect 202528 219218 202570 219454
rect 202806 219218 202848 219454
rect 202528 219134 202848 219218
rect 202528 218898 202570 219134
rect 202806 218898 202848 219134
rect 202528 218866 202848 218898
rect 233248 219454 233568 219486
rect 233248 219218 233290 219454
rect 233526 219218 233568 219454
rect 233248 219134 233568 219218
rect 233248 218898 233290 219134
rect 233526 218898 233568 219134
rect 233248 218866 233568 218898
rect 263968 219454 264288 219486
rect 263968 219218 264010 219454
rect 264246 219218 264288 219454
rect 263968 219134 264288 219218
rect 263968 218898 264010 219134
rect 264246 218898 264288 219134
rect 263968 218866 264288 218898
rect 294688 219454 295008 219486
rect 294688 219218 294730 219454
rect 294966 219218 295008 219454
rect 294688 219134 295008 219218
rect 294688 218898 294730 219134
rect 294966 218898 295008 219134
rect 294688 218866 295008 218898
rect 325408 219454 325728 219486
rect 325408 219218 325450 219454
rect 325686 219218 325728 219454
rect 325408 219134 325728 219218
rect 325408 218898 325450 219134
rect 325686 218898 325728 219134
rect 325408 218866 325728 218898
rect 356128 219454 356448 219486
rect 356128 219218 356170 219454
rect 356406 219218 356448 219454
rect 356128 219134 356448 219218
rect 356128 218898 356170 219134
rect 356406 218898 356448 219134
rect 356128 218866 356448 218898
rect 386848 219454 387168 219486
rect 386848 219218 386890 219454
rect 387126 219218 387168 219454
rect 386848 219134 387168 219218
rect 386848 218898 386890 219134
rect 387126 218898 387168 219134
rect 386848 218866 387168 218898
rect 417568 219454 417888 219486
rect 417568 219218 417610 219454
rect 417846 219218 417888 219454
rect 417568 219134 417888 219218
rect 417568 218898 417610 219134
rect 417846 218898 417888 219134
rect 417568 218866 417888 218898
rect 448288 219454 448608 219486
rect 448288 219218 448330 219454
rect 448566 219218 448608 219454
rect 448288 219134 448608 219218
rect 448288 218898 448330 219134
rect 448566 218898 448608 219134
rect 448288 218866 448608 218898
rect 479008 219454 479328 219486
rect 479008 219218 479050 219454
rect 479286 219218 479328 219454
rect 479008 219134 479328 219218
rect 479008 218898 479050 219134
rect 479286 218898 479328 219134
rect 479008 218866 479328 218898
rect 509728 219454 510048 219486
rect 509728 219218 509770 219454
rect 510006 219218 510048 219454
rect 509728 219134 510048 219218
rect 509728 218898 509770 219134
rect 510006 218898 510048 219134
rect 509728 218866 510048 218898
rect 540448 219454 540768 219486
rect 540448 219218 540490 219454
rect 540726 219218 540768 219454
rect 540448 219134 540768 219218
rect 540448 218898 540490 219134
rect 540726 218898 540768 219134
rect 540448 218866 540768 218898
rect 33568 201454 33888 201486
rect 33568 201218 33610 201454
rect 33846 201218 33888 201454
rect 33568 201134 33888 201218
rect 33568 200898 33610 201134
rect 33846 200898 33888 201134
rect 33568 200866 33888 200898
rect 64288 201454 64608 201486
rect 64288 201218 64330 201454
rect 64566 201218 64608 201454
rect 64288 201134 64608 201218
rect 64288 200898 64330 201134
rect 64566 200898 64608 201134
rect 64288 200866 64608 200898
rect 95008 201454 95328 201486
rect 95008 201218 95050 201454
rect 95286 201218 95328 201454
rect 95008 201134 95328 201218
rect 95008 200898 95050 201134
rect 95286 200898 95328 201134
rect 95008 200866 95328 200898
rect 125728 201454 126048 201486
rect 125728 201218 125770 201454
rect 126006 201218 126048 201454
rect 125728 201134 126048 201218
rect 125728 200898 125770 201134
rect 126006 200898 126048 201134
rect 125728 200866 126048 200898
rect 156448 201454 156768 201486
rect 156448 201218 156490 201454
rect 156726 201218 156768 201454
rect 156448 201134 156768 201218
rect 156448 200898 156490 201134
rect 156726 200898 156768 201134
rect 156448 200866 156768 200898
rect 187168 201454 187488 201486
rect 187168 201218 187210 201454
rect 187446 201218 187488 201454
rect 187168 201134 187488 201218
rect 187168 200898 187210 201134
rect 187446 200898 187488 201134
rect 187168 200866 187488 200898
rect 217888 201454 218208 201486
rect 217888 201218 217930 201454
rect 218166 201218 218208 201454
rect 217888 201134 218208 201218
rect 217888 200898 217930 201134
rect 218166 200898 218208 201134
rect 217888 200866 218208 200898
rect 248608 201454 248928 201486
rect 248608 201218 248650 201454
rect 248886 201218 248928 201454
rect 248608 201134 248928 201218
rect 248608 200898 248650 201134
rect 248886 200898 248928 201134
rect 248608 200866 248928 200898
rect 279328 201454 279648 201486
rect 279328 201218 279370 201454
rect 279606 201218 279648 201454
rect 279328 201134 279648 201218
rect 279328 200898 279370 201134
rect 279606 200898 279648 201134
rect 279328 200866 279648 200898
rect 310048 201454 310368 201486
rect 310048 201218 310090 201454
rect 310326 201218 310368 201454
rect 310048 201134 310368 201218
rect 310048 200898 310090 201134
rect 310326 200898 310368 201134
rect 310048 200866 310368 200898
rect 340768 201454 341088 201486
rect 340768 201218 340810 201454
rect 341046 201218 341088 201454
rect 340768 201134 341088 201218
rect 340768 200898 340810 201134
rect 341046 200898 341088 201134
rect 340768 200866 341088 200898
rect 371488 201454 371808 201486
rect 371488 201218 371530 201454
rect 371766 201218 371808 201454
rect 371488 201134 371808 201218
rect 371488 200898 371530 201134
rect 371766 200898 371808 201134
rect 371488 200866 371808 200898
rect 402208 201454 402528 201486
rect 402208 201218 402250 201454
rect 402486 201218 402528 201454
rect 402208 201134 402528 201218
rect 402208 200898 402250 201134
rect 402486 200898 402528 201134
rect 402208 200866 402528 200898
rect 432928 201454 433248 201486
rect 432928 201218 432970 201454
rect 433206 201218 433248 201454
rect 432928 201134 433248 201218
rect 432928 200898 432970 201134
rect 433206 200898 433248 201134
rect 432928 200866 433248 200898
rect 463648 201454 463968 201486
rect 463648 201218 463690 201454
rect 463926 201218 463968 201454
rect 463648 201134 463968 201218
rect 463648 200898 463690 201134
rect 463926 200898 463968 201134
rect 463648 200866 463968 200898
rect 494368 201454 494688 201486
rect 494368 201218 494410 201454
rect 494646 201218 494688 201454
rect 494368 201134 494688 201218
rect 494368 200898 494410 201134
rect 494646 200898 494688 201134
rect 494368 200866 494688 200898
rect 525088 201454 525408 201486
rect 525088 201218 525130 201454
rect 525366 201218 525408 201454
rect 525088 201134 525408 201218
rect 525088 200898 525130 201134
rect 525366 200898 525408 201134
rect 525088 200866 525408 200898
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 18208 183454 18528 183486
rect 18208 183218 18250 183454
rect 18486 183218 18528 183454
rect 18208 183134 18528 183218
rect 18208 182898 18250 183134
rect 18486 182898 18528 183134
rect 18208 182866 18528 182898
rect 48928 183454 49248 183486
rect 48928 183218 48970 183454
rect 49206 183218 49248 183454
rect 48928 183134 49248 183218
rect 48928 182898 48970 183134
rect 49206 182898 49248 183134
rect 48928 182866 49248 182898
rect 79648 183454 79968 183486
rect 79648 183218 79690 183454
rect 79926 183218 79968 183454
rect 79648 183134 79968 183218
rect 79648 182898 79690 183134
rect 79926 182898 79968 183134
rect 79648 182866 79968 182898
rect 110368 183454 110688 183486
rect 110368 183218 110410 183454
rect 110646 183218 110688 183454
rect 110368 183134 110688 183218
rect 110368 182898 110410 183134
rect 110646 182898 110688 183134
rect 110368 182866 110688 182898
rect 141088 183454 141408 183486
rect 141088 183218 141130 183454
rect 141366 183218 141408 183454
rect 141088 183134 141408 183218
rect 141088 182898 141130 183134
rect 141366 182898 141408 183134
rect 141088 182866 141408 182898
rect 171808 183454 172128 183486
rect 171808 183218 171850 183454
rect 172086 183218 172128 183454
rect 171808 183134 172128 183218
rect 171808 182898 171850 183134
rect 172086 182898 172128 183134
rect 171808 182866 172128 182898
rect 202528 183454 202848 183486
rect 202528 183218 202570 183454
rect 202806 183218 202848 183454
rect 202528 183134 202848 183218
rect 202528 182898 202570 183134
rect 202806 182898 202848 183134
rect 202528 182866 202848 182898
rect 233248 183454 233568 183486
rect 233248 183218 233290 183454
rect 233526 183218 233568 183454
rect 233248 183134 233568 183218
rect 233248 182898 233290 183134
rect 233526 182898 233568 183134
rect 233248 182866 233568 182898
rect 263968 183454 264288 183486
rect 263968 183218 264010 183454
rect 264246 183218 264288 183454
rect 263968 183134 264288 183218
rect 263968 182898 264010 183134
rect 264246 182898 264288 183134
rect 263968 182866 264288 182898
rect 294688 183454 295008 183486
rect 294688 183218 294730 183454
rect 294966 183218 295008 183454
rect 294688 183134 295008 183218
rect 294688 182898 294730 183134
rect 294966 182898 295008 183134
rect 294688 182866 295008 182898
rect 325408 183454 325728 183486
rect 325408 183218 325450 183454
rect 325686 183218 325728 183454
rect 325408 183134 325728 183218
rect 325408 182898 325450 183134
rect 325686 182898 325728 183134
rect 325408 182866 325728 182898
rect 356128 183454 356448 183486
rect 356128 183218 356170 183454
rect 356406 183218 356448 183454
rect 356128 183134 356448 183218
rect 356128 182898 356170 183134
rect 356406 182898 356448 183134
rect 356128 182866 356448 182898
rect 386848 183454 387168 183486
rect 386848 183218 386890 183454
rect 387126 183218 387168 183454
rect 386848 183134 387168 183218
rect 386848 182898 386890 183134
rect 387126 182898 387168 183134
rect 386848 182866 387168 182898
rect 417568 183454 417888 183486
rect 417568 183218 417610 183454
rect 417846 183218 417888 183454
rect 417568 183134 417888 183218
rect 417568 182898 417610 183134
rect 417846 182898 417888 183134
rect 417568 182866 417888 182898
rect 448288 183454 448608 183486
rect 448288 183218 448330 183454
rect 448566 183218 448608 183454
rect 448288 183134 448608 183218
rect 448288 182898 448330 183134
rect 448566 182898 448608 183134
rect 448288 182866 448608 182898
rect 479008 183454 479328 183486
rect 479008 183218 479050 183454
rect 479286 183218 479328 183454
rect 479008 183134 479328 183218
rect 479008 182898 479050 183134
rect 479286 182898 479328 183134
rect 479008 182866 479328 182898
rect 509728 183454 510048 183486
rect 509728 183218 509770 183454
rect 510006 183218 510048 183454
rect 509728 183134 510048 183218
rect 509728 182898 509770 183134
rect 510006 182898 510048 183134
rect 509728 182866 510048 182898
rect 540448 183454 540768 183486
rect 540448 183218 540490 183454
rect 540726 183218 540768 183454
rect 540448 183134 540768 183218
rect 540448 182898 540490 183134
rect 540726 182898 540768 183134
rect 540448 182866 540768 182898
rect 33568 165454 33888 165486
rect 33568 165218 33610 165454
rect 33846 165218 33888 165454
rect 33568 165134 33888 165218
rect 33568 164898 33610 165134
rect 33846 164898 33888 165134
rect 33568 164866 33888 164898
rect 64288 165454 64608 165486
rect 64288 165218 64330 165454
rect 64566 165218 64608 165454
rect 64288 165134 64608 165218
rect 64288 164898 64330 165134
rect 64566 164898 64608 165134
rect 64288 164866 64608 164898
rect 95008 165454 95328 165486
rect 95008 165218 95050 165454
rect 95286 165218 95328 165454
rect 95008 165134 95328 165218
rect 95008 164898 95050 165134
rect 95286 164898 95328 165134
rect 95008 164866 95328 164898
rect 125728 165454 126048 165486
rect 125728 165218 125770 165454
rect 126006 165218 126048 165454
rect 125728 165134 126048 165218
rect 125728 164898 125770 165134
rect 126006 164898 126048 165134
rect 125728 164866 126048 164898
rect 156448 165454 156768 165486
rect 156448 165218 156490 165454
rect 156726 165218 156768 165454
rect 156448 165134 156768 165218
rect 156448 164898 156490 165134
rect 156726 164898 156768 165134
rect 156448 164866 156768 164898
rect 187168 165454 187488 165486
rect 187168 165218 187210 165454
rect 187446 165218 187488 165454
rect 187168 165134 187488 165218
rect 187168 164898 187210 165134
rect 187446 164898 187488 165134
rect 187168 164866 187488 164898
rect 217888 165454 218208 165486
rect 217888 165218 217930 165454
rect 218166 165218 218208 165454
rect 217888 165134 218208 165218
rect 217888 164898 217930 165134
rect 218166 164898 218208 165134
rect 217888 164866 218208 164898
rect 248608 165454 248928 165486
rect 248608 165218 248650 165454
rect 248886 165218 248928 165454
rect 248608 165134 248928 165218
rect 248608 164898 248650 165134
rect 248886 164898 248928 165134
rect 248608 164866 248928 164898
rect 279328 165454 279648 165486
rect 279328 165218 279370 165454
rect 279606 165218 279648 165454
rect 279328 165134 279648 165218
rect 279328 164898 279370 165134
rect 279606 164898 279648 165134
rect 279328 164866 279648 164898
rect 310048 165454 310368 165486
rect 310048 165218 310090 165454
rect 310326 165218 310368 165454
rect 310048 165134 310368 165218
rect 310048 164898 310090 165134
rect 310326 164898 310368 165134
rect 310048 164866 310368 164898
rect 340768 165454 341088 165486
rect 340768 165218 340810 165454
rect 341046 165218 341088 165454
rect 340768 165134 341088 165218
rect 340768 164898 340810 165134
rect 341046 164898 341088 165134
rect 340768 164866 341088 164898
rect 371488 165454 371808 165486
rect 371488 165218 371530 165454
rect 371766 165218 371808 165454
rect 371488 165134 371808 165218
rect 371488 164898 371530 165134
rect 371766 164898 371808 165134
rect 371488 164866 371808 164898
rect 402208 165454 402528 165486
rect 402208 165218 402250 165454
rect 402486 165218 402528 165454
rect 402208 165134 402528 165218
rect 402208 164898 402250 165134
rect 402486 164898 402528 165134
rect 402208 164866 402528 164898
rect 432928 165454 433248 165486
rect 432928 165218 432970 165454
rect 433206 165218 433248 165454
rect 432928 165134 433248 165218
rect 432928 164898 432970 165134
rect 433206 164898 433248 165134
rect 432928 164866 433248 164898
rect 463648 165454 463968 165486
rect 463648 165218 463690 165454
rect 463926 165218 463968 165454
rect 463648 165134 463968 165218
rect 463648 164898 463690 165134
rect 463926 164898 463968 165134
rect 463648 164866 463968 164898
rect 494368 165454 494688 165486
rect 494368 165218 494410 165454
rect 494646 165218 494688 165454
rect 494368 165134 494688 165218
rect 494368 164898 494410 165134
rect 494646 164898 494688 165134
rect 494368 164866 494688 164898
rect 525088 165454 525408 165486
rect 525088 165218 525130 165454
rect 525366 165218 525408 165454
rect 525088 165134 525408 165218
rect 525088 164898 525130 165134
rect 525366 164898 525408 165134
rect 525088 164866 525408 164898
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 18208 147454 18528 147486
rect 18208 147218 18250 147454
rect 18486 147218 18528 147454
rect 18208 147134 18528 147218
rect 18208 146898 18250 147134
rect 18486 146898 18528 147134
rect 18208 146866 18528 146898
rect 48928 147454 49248 147486
rect 48928 147218 48970 147454
rect 49206 147218 49248 147454
rect 48928 147134 49248 147218
rect 48928 146898 48970 147134
rect 49206 146898 49248 147134
rect 48928 146866 49248 146898
rect 79648 147454 79968 147486
rect 79648 147218 79690 147454
rect 79926 147218 79968 147454
rect 79648 147134 79968 147218
rect 79648 146898 79690 147134
rect 79926 146898 79968 147134
rect 79648 146866 79968 146898
rect 110368 147454 110688 147486
rect 110368 147218 110410 147454
rect 110646 147218 110688 147454
rect 110368 147134 110688 147218
rect 110368 146898 110410 147134
rect 110646 146898 110688 147134
rect 110368 146866 110688 146898
rect 141088 147454 141408 147486
rect 141088 147218 141130 147454
rect 141366 147218 141408 147454
rect 141088 147134 141408 147218
rect 141088 146898 141130 147134
rect 141366 146898 141408 147134
rect 141088 146866 141408 146898
rect 171808 147454 172128 147486
rect 171808 147218 171850 147454
rect 172086 147218 172128 147454
rect 171808 147134 172128 147218
rect 171808 146898 171850 147134
rect 172086 146898 172128 147134
rect 171808 146866 172128 146898
rect 202528 147454 202848 147486
rect 202528 147218 202570 147454
rect 202806 147218 202848 147454
rect 202528 147134 202848 147218
rect 202528 146898 202570 147134
rect 202806 146898 202848 147134
rect 202528 146866 202848 146898
rect 233248 147454 233568 147486
rect 233248 147218 233290 147454
rect 233526 147218 233568 147454
rect 233248 147134 233568 147218
rect 233248 146898 233290 147134
rect 233526 146898 233568 147134
rect 233248 146866 233568 146898
rect 263968 147454 264288 147486
rect 263968 147218 264010 147454
rect 264246 147218 264288 147454
rect 263968 147134 264288 147218
rect 263968 146898 264010 147134
rect 264246 146898 264288 147134
rect 263968 146866 264288 146898
rect 294688 147454 295008 147486
rect 294688 147218 294730 147454
rect 294966 147218 295008 147454
rect 294688 147134 295008 147218
rect 294688 146898 294730 147134
rect 294966 146898 295008 147134
rect 294688 146866 295008 146898
rect 325408 147454 325728 147486
rect 325408 147218 325450 147454
rect 325686 147218 325728 147454
rect 325408 147134 325728 147218
rect 325408 146898 325450 147134
rect 325686 146898 325728 147134
rect 325408 146866 325728 146898
rect 356128 147454 356448 147486
rect 356128 147218 356170 147454
rect 356406 147218 356448 147454
rect 356128 147134 356448 147218
rect 356128 146898 356170 147134
rect 356406 146898 356448 147134
rect 356128 146866 356448 146898
rect 386848 147454 387168 147486
rect 386848 147218 386890 147454
rect 387126 147218 387168 147454
rect 386848 147134 387168 147218
rect 386848 146898 386890 147134
rect 387126 146898 387168 147134
rect 386848 146866 387168 146898
rect 417568 147454 417888 147486
rect 417568 147218 417610 147454
rect 417846 147218 417888 147454
rect 417568 147134 417888 147218
rect 417568 146898 417610 147134
rect 417846 146898 417888 147134
rect 417568 146866 417888 146898
rect 448288 147454 448608 147486
rect 448288 147218 448330 147454
rect 448566 147218 448608 147454
rect 448288 147134 448608 147218
rect 448288 146898 448330 147134
rect 448566 146898 448608 147134
rect 448288 146866 448608 146898
rect 479008 147454 479328 147486
rect 479008 147218 479050 147454
rect 479286 147218 479328 147454
rect 479008 147134 479328 147218
rect 479008 146898 479050 147134
rect 479286 146898 479328 147134
rect 479008 146866 479328 146898
rect 509728 147454 510048 147486
rect 509728 147218 509770 147454
rect 510006 147218 510048 147454
rect 509728 147134 510048 147218
rect 509728 146898 509770 147134
rect 510006 146898 510048 147134
rect 509728 146866 510048 146898
rect 540448 147454 540768 147486
rect 540448 147218 540490 147454
rect 540726 147218 540768 147454
rect 540448 147134 540768 147218
rect 540448 146898 540490 147134
rect 540726 146898 540768 147134
rect 540448 146866 540768 146898
rect 33568 129454 33888 129486
rect 33568 129218 33610 129454
rect 33846 129218 33888 129454
rect 33568 129134 33888 129218
rect 33568 128898 33610 129134
rect 33846 128898 33888 129134
rect 33568 128866 33888 128898
rect 64288 129454 64608 129486
rect 64288 129218 64330 129454
rect 64566 129218 64608 129454
rect 64288 129134 64608 129218
rect 64288 128898 64330 129134
rect 64566 128898 64608 129134
rect 64288 128866 64608 128898
rect 95008 129454 95328 129486
rect 95008 129218 95050 129454
rect 95286 129218 95328 129454
rect 95008 129134 95328 129218
rect 95008 128898 95050 129134
rect 95286 128898 95328 129134
rect 95008 128866 95328 128898
rect 125728 129454 126048 129486
rect 125728 129218 125770 129454
rect 126006 129218 126048 129454
rect 125728 129134 126048 129218
rect 125728 128898 125770 129134
rect 126006 128898 126048 129134
rect 125728 128866 126048 128898
rect 156448 129454 156768 129486
rect 156448 129218 156490 129454
rect 156726 129218 156768 129454
rect 156448 129134 156768 129218
rect 156448 128898 156490 129134
rect 156726 128898 156768 129134
rect 156448 128866 156768 128898
rect 187168 129454 187488 129486
rect 187168 129218 187210 129454
rect 187446 129218 187488 129454
rect 187168 129134 187488 129218
rect 187168 128898 187210 129134
rect 187446 128898 187488 129134
rect 187168 128866 187488 128898
rect 217888 129454 218208 129486
rect 217888 129218 217930 129454
rect 218166 129218 218208 129454
rect 217888 129134 218208 129218
rect 217888 128898 217930 129134
rect 218166 128898 218208 129134
rect 217888 128866 218208 128898
rect 248608 129454 248928 129486
rect 248608 129218 248650 129454
rect 248886 129218 248928 129454
rect 248608 129134 248928 129218
rect 248608 128898 248650 129134
rect 248886 128898 248928 129134
rect 248608 128866 248928 128898
rect 279328 129454 279648 129486
rect 279328 129218 279370 129454
rect 279606 129218 279648 129454
rect 279328 129134 279648 129218
rect 279328 128898 279370 129134
rect 279606 128898 279648 129134
rect 279328 128866 279648 128898
rect 310048 129454 310368 129486
rect 310048 129218 310090 129454
rect 310326 129218 310368 129454
rect 310048 129134 310368 129218
rect 310048 128898 310090 129134
rect 310326 128898 310368 129134
rect 310048 128866 310368 128898
rect 340768 129454 341088 129486
rect 340768 129218 340810 129454
rect 341046 129218 341088 129454
rect 340768 129134 341088 129218
rect 340768 128898 340810 129134
rect 341046 128898 341088 129134
rect 340768 128866 341088 128898
rect 371488 129454 371808 129486
rect 371488 129218 371530 129454
rect 371766 129218 371808 129454
rect 371488 129134 371808 129218
rect 371488 128898 371530 129134
rect 371766 128898 371808 129134
rect 371488 128866 371808 128898
rect 402208 129454 402528 129486
rect 402208 129218 402250 129454
rect 402486 129218 402528 129454
rect 402208 129134 402528 129218
rect 402208 128898 402250 129134
rect 402486 128898 402528 129134
rect 402208 128866 402528 128898
rect 432928 129454 433248 129486
rect 432928 129218 432970 129454
rect 433206 129218 433248 129454
rect 432928 129134 433248 129218
rect 432928 128898 432970 129134
rect 433206 128898 433248 129134
rect 432928 128866 433248 128898
rect 463648 129454 463968 129486
rect 463648 129218 463690 129454
rect 463926 129218 463968 129454
rect 463648 129134 463968 129218
rect 463648 128898 463690 129134
rect 463926 128898 463968 129134
rect 463648 128866 463968 128898
rect 494368 129454 494688 129486
rect 494368 129218 494410 129454
rect 494646 129218 494688 129454
rect 494368 129134 494688 129218
rect 494368 128898 494410 129134
rect 494646 128898 494688 129134
rect 494368 128866 494688 128898
rect 525088 129454 525408 129486
rect 525088 129218 525130 129454
rect 525366 129218 525408 129454
rect 525088 129134 525408 129218
rect 525088 128898 525130 129134
rect 525366 128898 525408 129134
rect 525088 128866 525408 128898
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 18208 111454 18528 111486
rect 18208 111218 18250 111454
rect 18486 111218 18528 111454
rect 18208 111134 18528 111218
rect 18208 110898 18250 111134
rect 18486 110898 18528 111134
rect 18208 110866 18528 110898
rect 48928 111454 49248 111486
rect 48928 111218 48970 111454
rect 49206 111218 49248 111454
rect 48928 111134 49248 111218
rect 48928 110898 48970 111134
rect 49206 110898 49248 111134
rect 48928 110866 49248 110898
rect 79648 111454 79968 111486
rect 79648 111218 79690 111454
rect 79926 111218 79968 111454
rect 79648 111134 79968 111218
rect 79648 110898 79690 111134
rect 79926 110898 79968 111134
rect 79648 110866 79968 110898
rect 110368 111454 110688 111486
rect 110368 111218 110410 111454
rect 110646 111218 110688 111454
rect 110368 111134 110688 111218
rect 110368 110898 110410 111134
rect 110646 110898 110688 111134
rect 110368 110866 110688 110898
rect 141088 111454 141408 111486
rect 141088 111218 141130 111454
rect 141366 111218 141408 111454
rect 141088 111134 141408 111218
rect 141088 110898 141130 111134
rect 141366 110898 141408 111134
rect 141088 110866 141408 110898
rect 171808 111454 172128 111486
rect 171808 111218 171850 111454
rect 172086 111218 172128 111454
rect 171808 111134 172128 111218
rect 171808 110898 171850 111134
rect 172086 110898 172128 111134
rect 171808 110866 172128 110898
rect 202528 111454 202848 111486
rect 202528 111218 202570 111454
rect 202806 111218 202848 111454
rect 202528 111134 202848 111218
rect 202528 110898 202570 111134
rect 202806 110898 202848 111134
rect 202528 110866 202848 110898
rect 233248 111454 233568 111486
rect 233248 111218 233290 111454
rect 233526 111218 233568 111454
rect 233248 111134 233568 111218
rect 233248 110898 233290 111134
rect 233526 110898 233568 111134
rect 233248 110866 233568 110898
rect 263968 111454 264288 111486
rect 263968 111218 264010 111454
rect 264246 111218 264288 111454
rect 263968 111134 264288 111218
rect 263968 110898 264010 111134
rect 264246 110898 264288 111134
rect 263968 110866 264288 110898
rect 294688 111454 295008 111486
rect 294688 111218 294730 111454
rect 294966 111218 295008 111454
rect 294688 111134 295008 111218
rect 294688 110898 294730 111134
rect 294966 110898 295008 111134
rect 294688 110866 295008 110898
rect 325408 111454 325728 111486
rect 325408 111218 325450 111454
rect 325686 111218 325728 111454
rect 325408 111134 325728 111218
rect 325408 110898 325450 111134
rect 325686 110898 325728 111134
rect 325408 110866 325728 110898
rect 356128 111454 356448 111486
rect 356128 111218 356170 111454
rect 356406 111218 356448 111454
rect 356128 111134 356448 111218
rect 356128 110898 356170 111134
rect 356406 110898 356448 111134
rect 356128 110866 356448 110898
rect 386848 111454 387168 111486
rect 386848 111218 386890 111454
rect 387126 111218 387168 111454
rect 386848 111134 387168 111218
rect 386848 110898 386890 111134
rect 387126 110898 387168 111134
rect 386848 110866 387168 110898
rect 417568 111454 417888 111486
rect 417568 111218 417610 111454
rect 417846 111218 417888 111454
rect 417568 111134 417888 111218
rect 417568 110898 417610 111134
rect 417846 110898 417888 111134
rect 417568 110866 417888 110898
rect 448288 111454 448608 111486
rect 448288 111218 448330 111454
rect 448566 111218 448608 111454
rect 448288 111134 448608 111218
rect 448288 110898 448330 111134
rect 448566 110898 448608 111134
rect 448288 110866 448608 110898
rect 479008 111454 479328 111486
rect 479008 111218 479050 111454
rect 479286 111218 479328 111454
rect 479008 111134 479328 111218
rect 479008 110898 479050 111134
rect 479286 110898 479328 111134
rect 479008 110866 479328 110898
rect 509728 111454 510048 111486
rect 509728 111218 509770 111454
rect 510006 111218 510048 111454
rect 509728 111134 510048 111218
rect 509728 110898 509770 111134
rect 510006 110898 510048 111134
rect 509728 110866 510048 110898
rect 540448 111454 540768 111486
rect 540448 111218 540490 111454
rect 540726 111218 540768 111454
rect 540448 111134 540768 111218
rect 540448 110898 540490 111134
rect 540726 110898 540768 111134
rect 540448 110866 540768 110898
rect 33568 93454 33888 93486
rect 33568 93218 33610 93454
rect 33846 93218 33888 93454
rect 33568 93134 33888 93218
rect 33568 92898 33610 93134
rect 33846 92898 33888 93134
rect 33568 92866 33888 92898
rect 64288 93454 64608 93486
rect 64288 93218 64330 93454
rect 64566 93218 64608 93454
rect 64288 93134 64608 93218
rect 64288 92898 64330 93134
rect 64566 92898 64608 93134
rect 64288 92866 64608 92898
rect 95008 93454 95328 93486
rect 95008 93218 95050 93454
rect 95286 93218 95328 93454
rect 95008 93134 95328 93218
rect 95008 92898 95050 93134
rect 95286 92898 95328 93134
rect 95008 92866 95328 92898
rect 125728 93454 126048 93486
rect 125728 93218 125770 93454
rect 126006 93218 126048 93454
rect 125728 93134 126048 93218
rect 125728 92898 125770 93134
rect 126006 92898 126048 93134
rect 125728 92866 126048 92898
rect 156448 93454 156768 93486
rect 156448 93218 156490 93454
rect 156726 93218 156768 93454
rect 156448 93134 156768 93218
rect 156448 92898 156490 93134
rect 156726 92898 156768 93134
rect 156448 92866 156768 92898
rect 187168 93454 187488 93486
rect 187168 93218 187210 93454
rect 187446 93218 187488 93454
rect 187168 93134 187488 93218
rect 187168 92898 187210 93134
rect 187446 92898 187488 93134
rect 187168 92866 187488 92898
rect 217888 93454 218208 93486
rect 217888 93218 217930 93454
rect 218166 93218 218208 93454
rect 217888 93134 218208 93218
rect 217888 92898 217930 93134
rect 218166 92898 218208 93134
rect 217888 92866 218208 92898
rect 248608 93454 248928 93486
rect 248608 93218 248650 93454
rect 248886 93218 248928 93454
rect 248608 93134 248928 93218
rect 248608 92898 248650 93134
rect 248886 92898 248928 93134
rect 248608 92866 248928 92898
rect 279328 93454 279648 93486
rect 279328 93218 279370 93454
rect 279606 93218 279648 93454
rect 279328 93134 279648 93218
rect 279328 92898 279370 93134
rect 279606 92898 279648 93134
rect 279328 92866 279648 92898
rect 310048 93454 310368 93486
rect 310048 93218 310090 93454
rect 310326 93218 310368 93454
rect 310048 93134 310368 93218
rect 310048 92898 310090 93134
rect 310326 92898 310368 93134
rect 310048 92866 310368 92898
rect 340768 93454 341088 93486
rect 340768 93218 340810 93454
rect 341046 93218 341088 93454
rect 340768 93134 341088 93218
rect 340768 92898 340810 93134
rect 341046 92898 341088 93134
rect 340768 92866 341088 92898
rect 371488 93454 371808 93486
rect 371488 93218 371530 93454
rect 371766 93218 371808 93454
rect 371488 93134 371808 93218
rect 371488 92898 371530 93134
rect 371766 92898 371808 93134
rect 371488 92866 371808 92898
rect 402208 93454 402528 93486
rect 402208 93218 402250 93454
rect 402486 93218 402528 93454
rect 402208 93134 402528 93218
rect 402208 92898 402250 93134
rect 402486 92898 402528 93134
rect 402208 92866 402528 92898
rect 432928 93454 433248 93486
rect 432928 93218 432970 93454
rect 433206 93218 433248 93454
rect 432928 93134 433248 93218
rect 432928 92898 432970 93134
rect 433206 92898 433248 93134
rect 432928 92866 433248 92898
rect 463648 93454 463968 93486
rect 463648 93218 463690 93454
rect 463926 93218 463968 93454
rect 463648 93134 463968 93218
rect 463648 92898 463690 93134
rect 463926 92898 463968 93134
rect 463648 92866 463968 92898
rect 494368 93454 494688 93486
rect 494368 93218 494410 93454
rect 494646 93218 494688 93454
rect 494368 93134 494688 93218
rect 494368 92898 494410 93134
rect 494646 92898 494688 93134
rect 494368 92866 494688 92898
rect 525088 93454 525408 93486
rect 525088 93218 525130 93454
rect 525366 93218 525408 93454
rect 525088 93134 525408 93218
rect 525088 92898 525130 93134
rect 525366 92898 525408 93134
rect 525088 92866 525408 92898
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 18208 75454 18528 75486
rect 18208 75218 18250 75454
rect 18486 75218 18528 75454
rect 18208 75134 18528 75218
rect 18208 74898 18250 75134
rect 18486 74898 18528 75134
rect 18208 74866 18528 74898
rect 48928 75454 49248 75486
rect 48928 75218 48970 75454
rect 49206 75218 49248 75454
rect 48928 75134 49248 75218
rect 48928 74898 48970 75134
rect 49206 74898 49248 75134
rect 48928 74866 49248 74898
rect 79648 75454 79968 75486
rect 79648 75218 79690 75454
rect 79926 75218 79968 75454
rect 79648 75134 79968 75218
rect 79648 74898 79690 75134
rect 79926 74898 79968 75134
rect 79648 74866 79968 74898
rect 110368 75454 110688 75486
rect 110368 75218 110410 75454
rect 110646 75218 110688 75454
rect 110368 75134 110688 75218
rect 110368 74898 110410 75134
rect 110646 74898 110688 75134
rect 110368 74866 110688 74898
rect 141088 75454 141408 75486
rect 141088 75218 141130 75454
rect 141366 75218 141408 75454
rect 141088 75134 141408 75218
rect 141088 74898 141130 75134
rect 141366 74898 141408 75134
rect 141088 74866 141408 74898
rect 171808 75454 172128 75486
rect 171808 75218 171850 75454
rect 172086 75218 172128 75454
rect 171808 75134 172128 75218
rect 171808 74898 171850 75134
rect 172086 74898 172128 75134
rect 171808 74866 172128 74898
rect 202528 75454 202848 75486
rect 202528 75218 202570 75454
rect 202806 75218 202848 75454
rect 202528 75134 202848 75218
rect 202528 74898 202570 75134
rect 202806 74898 202848 75134
rect 202528 74866 202848 74898
rect 233248 75454 233568 75486
rect 233248 75218 233290 75454
rect 233526 75218 233568 75454
rect 233248 75134 233568 75218
rect 233248 74898 233290 75134
rect 233526 74898 233568 75134
rect 233248 74866 233568 74898
rect 263968 75454 264288 75486
rect 263968 75218 264010 75454
rect 264246 75218 264288 75454
rect 263968 75134 264288 75218
rect 263968 74898 264010 75134
rect 264246 74898 264288 75134
rect 263968 74866 264288 74898
rect 294688 75454 295008 75486
rect 294688 75218 294730 75454
rect 294966 75218 295008 75454
rect 294688 75134 295008 75218
rect 294688 74898 294730 75134
rect 294966 74898 295008 75134
rect 294688 74866 295008 74898
rect 325408 75454 325728 75486
rect 325408 75218 325450 75454
rect 325686 75218 325728 75454
rect 325408 75134 325728 75218
rect 325408 74898 325450 75134
rect 325686 74898 325728 75134
rect 325408 74866 325728 74898
rect 356128 75454 356448 75486
rect 356128 75218 356170 75454
rect 356406 75218 356448 75454
rect 356128 75134 356448 75218
rect 356128 74898 356170 75134
rect 356406 74898 356448 75134
rect 356128 74866 356448 74898
rect 386848 75454 387168 75486
rect 386848 75218 386890 75454
rect 387126 75218 387168 75454
rect 386848 75134 387168 75218
rect 386848 74898 386890 75134
rect 387126 74898 387168 75134
rect 386848 74866 387168 74898
rect 417568 75454 417888 75486
rect 417568 75218 417610 75454
rect 417846 75218 417888 75454
rect 417568 75134 417888 75218
rect 417568 74898 417610 75134
rect 417846 74898 417888 75134
rect 417568 74866 417888 74898
rect 448288 75454 448608 75486
rect 448288 75218 448330 75454
rect 448566 75218 448608 75454
rect 448288 75134 448608 75218
rect 448288 74898 448330 75134
rect 448566 74898 448608 75134
rect 448288 74866 448608 74898
rect 479008 75454 479328 75486
rect 479008 75218 479050 75454
rect 479286 75218 479328 75454
rect 479008 75134 479328 75218
rect 479008 74898 479050 75134
rect 479286 74898 479328 75134
rect 479008 74866 479328 74898
rect 509728 75454 510048 75486
rect 509728 75218 509770 75454
rect 510006 75218 510048 75454
rect 509728 75134 510048 75218
rect 509728 74898 509770 75134
rect 510006 74898 510048 75134
rect 509728 74866 510048 74898
rect 540448 75454 540768 75486
rect 540448 75218 540490 75454
rect 540726 75218 540768 75454
rect 540448 75134 540768 75218
rect 540448 74898 540490 75134
rect 540726 74898 540768 75134
rect 540448 74866 540768 74898
rect 33568 57454 33888 57486
rect 33568 57218 33610 57454
rect 33846 57218 33888 57454
rect 33568 57134 33888 57218
rect 33568 56898 33610 57134
rect 33846 56898 33888 57134
rect 33568 56866 33888 56898
rect 64288 57454 64608 57486
rect 64288 57218 64330 57454
rect 64566 57218 64608 57454
rect 64288 57134 64608 57218
rect 64288 56898 64330 57134
rect 64566 56898 64608 57134
rect 64288 56866 64608 56898
rect 95008 57454 95328 57486
rect 95008 57218 95050 57454
rect 95286 57218 95328 57454
rect 95008 57134 95328 57218
rect 95008 56898 95050 57134
rect 95286 56898 95328 57134
rect 95008 56866 95328 56898
rect 125728 57454 126048 57486
rect 125728 57218 125770 57454
rect 126006 57218 126048 57454
rect 125728 57134 126048 57218
rect 125728 56898 125770 57134
rect 126006 56898 126048 57134
rect 125728 56866 126048 56898
rect 156448 57454 156768 57486
rect 156448 57218 156490 57454
rect 156726 57218 156768 57454
rect 156448 57134 156768 57218
rect 156448 56898 156490 57134
rect 156726 56898 156768 57134
rect 156448 56866 156768 56898
rect 187168 57454 187488 57486
rect 187168 57218 187210 57454
rect 187446 57218 187488 57454
rect 187168 57134 187488 57218
rect 187168 56898 187210 57134
rect 187446 56898 187488 57134
rect 187168 56866 187488 56898
rect 217888 57454 218208 57486
rect 217888 57218 217930 57454
rect 218166 57218 218208 57454
rect 217888 57134 218208 57218
rect 217888 56898 217930 57134
rect 218166 56898 218208 57134
rect 217888 56866 218208 56898
rect 248608 57454 248928 57486
rect 248608 57218 248650 57454
rect 248886 57218 248928 57454
rect 248608 57134 248928 57218
rect 248608 56898 248650 57134
rect 248886 56898 248928 57134
rect 248608 56866 248928 56898
rect 279328 57454 279648 57486
rect 279328 57218 279370 57454
rect 279606 57218 279648 57454
rect 279328 57134 279648 57218
rect 279328 56898 279370 57134
rect 279606 56898 279648 57134
rect 279328 56866 279648 56898
rect 310048 57454 310368 57486
rect 310048 57218 310090 57454
rect 310326 57218 310368 57454
rect 310048 57134 310368 57218
rect 310048 56898 310090 57134
rect 310326 56898 310368 57134
rect 310048 56866 310368 56898
rect 340768 57454 341088 57486
rect 340768 57218 340810 57454
rect 341046 57218 341088 57454
rect 340768 57134 341088 57218
rect 340768 56898 340810 57134
rect 341046 56898 341088 57134
rect 340768 56866 341088 56898
rect 371488 57454 371808 57486
rect 371488 57218 371530 57454
rect 371766 57218 371808 57454
rect 371488 57134 371808 57218
rect 371488 56898 371530 57134
rect 371766 56898 371808 57134
rect 371488 56866 371808 56898
rect 402208 57454 402528 57486
rect 402208 57218 402250 57454
rect 402486 57218 402528 57454
rect 402208 57134 402528 57218
rect 402208 56898 402250 57134
rect 402486 56898 402528 57134
rect 402208 56866 402528 56898
rect 432928 57454 433248 57486
rect 432928 57218 432970 57454
rect 433206 57218 433248 57454
rect 432928 57134 433248 57218
rect 432928 56898 432970 57134
rect 433206 56898 433248 57134
rect 432928 56866 433248 56898
rect 463648 57454 463968 57486
rect 463648 57218 463690 57454
rect 463926 57218 463968 57454
rect 463648 57134 463968 57218
rect 463648 56898 463690 57134
rect 463926 56898 463968 57134
rect 463648 56866 463968 56898
rect 494368 57454 494688 57486
rect 494368 57218 494410 57454
rect 494646 57218 494688 57454
rect 494368 57134 494688 57218
rect 494368 56898 494410 57134
rect 494646 56898 494688 57134
rect 494368 56866 494688 56898
rect 525088 57454 525408 57486
rect 525088 57218 525130 57454
rect 525366 57218 525408 57454
rect 525088 57134 525408 57218
rect 525088 56898 525130 57134
rect 525366 56898 525408 57134
rect 525088 56866 525408 56898
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 14614 13574 48000
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 21454 20414 48000
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 25174 24134 48000
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 28894 27854 48000
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 32614 31574 48000
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 39454 38414 48000
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 43174 42134 48000
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 46894 45854 48000
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 48000
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 48000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 48000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 48000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 48000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 48000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 48000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 48000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 48000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 48000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 48000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 48000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 48000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 48000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 48000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 48000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 48000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 48000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 48000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 48000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 48000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 48000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 48000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 48000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 48000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 48000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 48000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 48000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 48000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 48000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 48000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 48000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 48000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 48000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 48000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 48000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 48000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 48000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 48000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 48000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 48000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 48000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 48000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 48000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 48000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 48000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 48000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 48000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 48000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 48000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 48000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 48000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 48000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 48000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 48000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 48000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 48000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 48000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 48000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 48000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 48000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 48000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 48000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 48000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 48000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 48000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 48000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 48000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 48000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 48000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 48000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 48000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 48000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 48000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 48000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 48000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 48000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 48000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 48000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 48000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 48000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 48000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 48000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 48000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 48000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 48000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 48000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 48000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 48000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 48000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 48000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 48000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 48000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 48000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 48000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 48000
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 48000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 48000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 48000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 48000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 48000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 48000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 48000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 48000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 48000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 48000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 48000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 28894 531854 48000
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 32614 535574 48000
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 39454 542414 48000
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 43174 546134 48000
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 46894 549854 48000
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 14614 553574 48000
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 18250 651218 18486 651454
rect 18250 650898 18486 651134
rect 48970 651218 49206 651454
rect 48970 650898 49206 651134
rect 79690 651218 79926 651454
rect 79690 650898 79926 651134
rect 110410 651218 110646 651454
rect 110410 650898 110646 651134
rect 141130 651218 141366 651454
rect 141130 650898 141366 651134
rect 171850 651218 172086 651454
rect 171850 650898 172086 651134
rect 202570 651218 202806 651454
rect 202570 650898 202806 651134
rect 233290 651218 233526 651454
rect 233290 650898 233526 651134
rect 264010 651218 264246 651454
rect 264010 650898 264246 651134
rect 294730 651218 294966 651454
rect 294730 650898 294966 651134
rect 325450 651218 325686 651454
rect 325450 650898 325686 651134
rect 356170 651218 356406 651454
rect 356170 650898 356406 651134
rect 386890 651218 387126 651454
rect 386890 650898 387126 651134
rect 417610 651218 417846 651454
rect 417610 650898 417846 651134
rect 448330 651218 448566 651454
rect 448330 650898 448566 651134
rect 479050 651218 479286 651454
rect 479050 650898 479286 651134
rect 509770 651218 510006 651454
rect 509770 650898 510006 651134
rect 540490 651218 540726 651454
rect 540490 650898 540726 651134
rect 33610 633218 33846 633454
rect 33610 632898 33846 633134
rect 64330 633218 64566 633454
rect 64330 632898 64566 633134
rect 95050 633218 95286 633454
rect 95050 632898 95286 633134
rect 125770 633218 126006 633454
rect 125770 632898 126006 633134
rect 156490 633218 156726 633454
rect 156490 632898 156726 633134
rect 187210 633218 187446 633454
rect 187210 632898 187446 633134
rect 217930 633218 218166 633454
rect 217930 632898 218166 633134
rect 248650 633218 248886 633454
rect 248650 632898 248886 633134
rect 279370 633218 279606 633454
rect 279370 632898 279606 633134
rect 310090 633218 310326 633454
rect 310090 632898 310326 633134
rect 340810 633218 341046 633454
rect 340810 632898 341046 633134
rect 371530 633218 371766 633454
rect 371530 632898 371766 633134
rect 402250 633218 402486 633454
rect 402250 632898 402486 633134
rect 432970 633218 433206 633454
rect 432970 632898 433206 633134
rect 463690 633218 463926 633454
rect 463690 632898 463926 633134
rect 494410 633218 494646 633454
rect 494410 632898 494646 633134
rect 525130 633218 525366 633454
rect 525130 632898 525366 633134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 18250 615218 18486 615454
rect 18250 614898 18486 615134
rect 48970 615218 49206 615454
rect 48970 614898 49206 615134
rect 79690 615218 79926 615454
rect 79690 614898 79926 615134
rect 110410 615218 110646 615454
rect 110410 614898 110646 615134
rect 141130 615218 141366 615454
rect 141130 614898 141366 615134
rect 171850 615218 172086 615454
rect 171850 614898 172086 615134
rect 202570 615218 202806 615454
rect 202570 614898 202806 615134
rect 233290 615218 233526 615454
rect 233290 614898 233526 615134
rect 264010 615218 264246 615454
rect 264010 614898 264246 615134
rect 294730 615218 294966 615454
rect 294730 614898 294966 615134
rect 325450 615218 325686 615454
rect 325450 614898 325686 615134
rect 356170 615218 356406 615454
rect 356170 614898 356406 615134
rect 386890 615218 387126 615454
rect 386890 614898 387126 615134
rect 417610 615218 417846 615454
rect 417610 614898 417846 615134
rect 448330 615218 448566 615454
rect 448330 614898 448566 615134
rect 479050 615218 479286 615454
rect 479050 614898 479286 615134
rect 509770 615218 510006 615454
rect 509770 614898 510006 615134
rect 540490 615218 540726 615454
rect 540490 614898 540726 615134
rect 33610 597218 33846 597454
rect 33610 596898 33846 597134
rect 64330 597218 64566 597454
rect 64330 596898 64566 597134
rect 95050 597218 95286 597454
rect 95050 596898 95286 597134
rect 125770 597218 126006 597454
rect 125770 596898 126006 597134
rect 156490 597218 156726 597454
rect 156490 596898 156726 597134
rect 187210 597218 187446 597454
rect 187210 596898 187446 597134
rect 217930 597218 218166 597454
rect 217930 596898 218166 597134
rect 248650 597218 248886 597454
rect 248650 596898 248886 597134
rect 279370 597218 279606 597454
rect 279370 596898 279606 597134
rect 310090 597218 310326 597454
rect 310090 596898 310326 597134
rect 340810 597218 341046 597454
rect 340810 596898 341046 597134
rect 371530 597218 371766 597454
rect 371530 596898 371766 597134
rect 402250 597218 402486 597454
rect 402250 596898 402486 597134
rect 432970 597218 433206 597454
rect 432970 596898 433206 597134
rect 463690 597218 463926 597454
rect 463690 596898 463926 597134
rect 494410 597218 494646 597454
rect 494410 596898 494646 597134
rect 525130 597218 525366 597454
rect 525130 596898 525366 597134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 18250 579218 18486 579454
rect 18250 578898 18486 579134
rect 48970 579218 49206 579454
rect 48970 578898 49206 579134
rect 79690 579218 79926 579454
rect 79690 578898 79926 579134
rect 110410 579218 110646 579454
rect 110410 578898 110646 579134
rect 141130 579218 141366 579454
rect 141130 578898 141366 579134
rect 171850 579218 172086 579454
rect 171850 578898 172086 579134
rect 202570 579218 202806 579454
rect 202570 578898 202806 579134
rect 233290 579218 233526 579454
rect 233290 578898 233526 579134
rect 264010 579218 264246 579454
rect 264010 578898 264246 579134
rect 294730 579218 294966 579454
rect 294730 578898 294966 579134
rect 325450 579218 325686 579454
rect 325450 578898 325686 579134
rect 356170 579218 356406 579454
rect 356170 578898 356406 579134
rect 386890 579218 387126 579454
rect 386890 578898 387126 579134
rect 417610 579218 417846 579454
rect 417610 578898 417846 579134
rect 448330 579218 448566 579454
rect 448330 578898 448566 579134
rect 479050 579218 479286 579454
rect 479050 578898 479286 579134
rect 509770 579218 510006 579454
rect 509770 578898 510006 579134
rect 540490 579218 540726 579454
rect 540490 578898 540726 579134
rect 33610 561218 33846 561454
rect 33610 560898 33846 561134
rect 64330 561218 64566 561454
rect 64330 560898 64566 561134
rect 95050 561218 95286 561454
rect 95050 560898 95286 561134
rect 125770 561218 126006 561454
rect 125770 560898 126006 561134
rect 156490 561218 156726 561454
rect 156490 560898 156726 561134
rect 187210 561218 187446 561454
rect 187210 560898 187446 561134
rect 217930 561218 218166 561454
rect 217930 560898 218166 561134
rect 248650 561218 248886 561454
rect 248650 560898 248886 561134
rect 279370 561218 279606 561454
rect 279370 560898 279606 561134
rect 310090 561218 310326 561454
rect 310090 560898 310326 561134
rect 340810 561218 341046 561454
rect 340810 560898 341046 561134
rect 371530 561218 371766 561454
rect 371530 560898 371766 561134
rect 402250 561218 402486 561454
rect 402250 560898 402486 561134
rect 432970 561218 433206 561454
rect 432970 560898 433206 561134
rect 463690 561218 463926 561454
rect 463690 560898 463926 561134
rect 494410 561218 494646 561454
rect 494410 560898 494646 561134
rect 525130 561218 525366 561454
rect 525130 560898 525366 561134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 18250 543218 18486 543454
rect 18250 542898 18486 543134
rect 48970 543218 49206 543454
rect 48970 542898 49206 543134
rect 79690 543218 79926 543454
rect 79690 542898 79926 543134
rect 110410 543218 110646 543454
rect 110410 542898 110646 543134
rect 141130 543218 141366 543454
rect 141130 542898 141366 543134
rect 171850 543218 172086 543454
rect 171850 542898 172086 543134
rect 202570 543218 202806 543454
rect 202570 542898 202806 543134
rect 233290 543218 233526 543454
rect 233290 542898 233526 543134
rect 264010 543218 264246 543454
rect 264010 542898 264246 543134
rect 294730 543218 294966 543454
rect 294730 542898 294966 543134
rect 325450 543218 325686 543454
rect 325450 542898 325686 543134
rect 356170 543218 356406 543454
rect 356170 542898 356406 543134
rect 386890 543218 387126 543454
rect 386890 542898 387126 543134
rect 417610 543218 417846 543454
rect 417610 542898 417846 543134
rect 448330 543218 448566 543454
rect 448330 542898 448566 543134
rect 479050 543218 479286 543454
rect 479050 542898 479286 543134
rect 509770 543218 510006 543454
rect 509770 542898 510006 543134
rect 540490 543218 540726 543454
rect 540490 542898 540726 543134
rect 33610 525218 33846 525454
rect 33610 524898 33846 525134
rect 64330 525218 64566 525454
rect 64330 524898 64566 525134
rect 95050 525218 95286 525454
rect 95050 524898 95286 525134
rect 125770 525218 126006 525454
rect 125770 524898 126006 525134
rect 156490 525218 156726 525454
rect 156490 524898 156726 525134
rect 187210 525218 187446 525454
rect 187210 524898 187446 525134
rect 217930 525218 218166 525454
rect 217930 524898 218166 525134
rect 248650 525218 248886 525454
rect 248650 524898 248886 525134
rect 279370 525218 279606 525454
rect 279370 524898 279606 525134
rect 310090 525218 310326 525454
rect 310090 524898 310326 525134
rect 340810 525218 341046 525454
rect 340810 524898 341046 525134
rect 371530 525218 371766 525454
rect 371530 524898 371766 525134
rect 402250 525218 402486 525454
rect 402250 524898 402486 525134
rect 432970 525218 433206 525454
rect 432970 524898 433206 525134
rect 463690 525218 463926 525454
rect 463690 524898 463926 525134
rect 494410 525218 494646 525454
rect 494410 524898 494646 525134
rect 525130 525218 525366 525454
rect 525130 524898 525366 525134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 18250 507218 18486 507454
rect 18250 506898 18486 507134
rect 48970 507218 49206 507454
rect 48970 506898 49206 507134
rect 79690 507218 79926 507454
rect 79690 506898 79926 507134
rect 110410 507218 110646 507454
rect 110410 506898 110646 507134
rect 141130 507218 141366 507454
rect 141130 506898 141366 507134
rect 171850 507218 172086 507454
rect 171850 506898 172086 507134
rect 202570 507218 202806 507454
rect 202570 506898 202806 507134
rect 233290 507218 233526 507454
rect 233290 506898 233526 507134
rect 264010 507218 264246 507454
rect 264010 506898 264246 507134
rect 294730 507218 294966 507454
rect 294730 506898 294966 507134
rect 325450 507218 325686 507454
rect 325450 506898 325686 507134
rect 356170 507218 356406 507454
rect 356170 506898 356406 507134
rect 386890 507218 387126 507454
rect 386890 506898 387126 507134
rect 417610 507218 417846 507454
rect 417610 506898 417846 507134
rect 448330 507218 448566 507454
rect 448330 506898 448566 507134
rect 479050 507218 479286 507454
rect 479050 506898 479286 507134
rect 509770 507218 510006 507454
rect 509770 506898 510006 507134
rect 540490 507218 540726 507454
rect 540490 506898 540726 507134
rect 33610 489218 33846 489454
rect 33610 488898 33846 489134
rect 64330 489218 64566 489454
rect 64330 488898 64566 489134
rect 95050 489218 95286 489454
rect 95050 488898 95286 489134
rect 125770 489218 126006 489454
rect 125770 488898 126006 489134
rect 156490 489218 156726 489454
rect 156490 488898 156726 489134
rect 187210 489218 187446 489454
rect 187210 488898 187446 489134
rect 217930 489218 218166 489454
rect 217930 488898 218166 489134
rect 248650 489218 248886 489454
rect 248650 488898 248886 489134
rect 279370 489218 279606 489454
rect 279370 488898 279606 489134
rect 310090 489218 310326 489454
rect 310090 488898 310326 489134
rect 340810 489218 341046 489454
rect 340810 488898 341046 489134
rect 371530 489218 371766 489454
rect 371530 488898 371766 489134
rect 402250 489218 402486 489454
rect 402250 488898 402486 489134
rect 432970 489218 433206 489454
rect 432970 488898 433206 489134
rect 463690 489218 463926 489454
rect 463690 488898 463926 489134
rect 494410 489218 494646 489454
rect 494410 488898 494646 489134
rect 525130 489218 525366 489454
rect 525130 488898 525366 489134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 18250 471218 18486 471454
rect 18250 470898 18486 471134
rect 48970 471218 49206 471454
rect 48970 470898 49206 471134
rect 79690 471218 79926 471454
rect 79690 470898 79926 471134
rect 110410 471218 110646 471454
rect 110410 470898 110646 471134
rect 141130 471218 141366 471454
rect 141130 470898 141366 471134
rect 171850 471218 172086 471454
rect 171850 470898 172086 471134
rect 202570 471218 202806 471454
rect 202570 470898 202806 471134
rect 233290 471218 233526 471454
rect 233290 470898 233526 471134
rect 264010 471218 264246 471454
rect 264010 470898 264246 471134
rect 294730 471218 294966 471454
rect 294730 470898 294966 471134
rect 325450 471218 325686 471454
rect 325450 470898 325686 471134
rect 356170 471218 356406 471454
rect 356170 470898 356406 471134
rect 386890 471218 387126 471454
rect 386890 470898 387126 471134
rect 417610 471218 417846 471454
rect 417610 470898 417846 471134
rect 448330 471218 448566 471454
rect 448330 470898 448566 471134
rect 479050 471218 479286 471454
rect 479050 470898 479286 471134
rect 509770 471218 510006 471454
rect 509770 470898 510006 471134
rect 540490 471218 540726 471454
rect 540490 470898 540726 471134
rect 33610 453218 33846 453454
rect 33610 452898 33846 453134
rect 64330 453218 64566 453454
rect 64330 452898 64566 453134
rect 95050 453218 95286 453454
rect 95050 452898 95286 453134
rect 125770 453218 126006 453454
rect 125770 452898 126006 453134
rect 156490 453218 156726 453454
rect 156490 452898 156726 453134
rect 187210 453218 187446 453454
rect 187210 452898 187446 453134
rect 217930 453218 218166 453454
rect 217930 452898 218166 453134
rect 248650 453218 248886 453454
rect 248650 452898 248886 453134
rect 279370 453218 279606 453454
rect 279370 452898 279606 453134
rect 310090 453218 310326 453454
rect 310090 452898 310326 453134
rect 340810 453218 341046 453454
rect 340810 452898 341046 453134
rect 371530 453218 371766 453454
rect 371530 452898 371766 453134
rect 402250 453218 402486 453454
rect 402250 452898 402486 453134
rect 432970 453218 433206 453454
rect 432970 452898 433206 453134
rect 463690 453218 463926 453454
rect 463690 452898 463926 453134
rect 494410 453218 494646 453454
rect 494410 452898 494646 453134
rect 525130 453218 525366 453454
rect 525130 452898 525366 453134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 18250 435218 18486 435454
rect 18250 434898 18486 435134
rect 48970 435218 49206 435454
rect 48970 434898 49206 435134
rect 79690 435218 79926 435454
rect 79690 434898 79926 435134
rect 110410 435218 110646 435454
rect 110410 434898 110646 435134
rect 141130 435218 141366 435454
rect 141130 434898 141366 435134
rect 171850 435218 172086 435454
rect 171850 434898 172086 435134
rect 202570 435218 202806 435454
rect 202570 434898 202806 435134
rect 233290 435218 233526 435454
rect 233290 434898 233526 435134
rect 264010 435218 264246 435454
rect 264010 434898 264246 435134
rect 294730 435218 294966 435454
rect 294730 434898 294966 435134
rect 325450 435218 325686 435454
rect 325450 434898 325686 435134
rect 356170 435218 356406 435454
rect 356170 434898 356406 435134
rect 386890 435218 387126 435454
rect 386890 434898 387126 435134
rect 417610 435218 417846 435454
rect 417610 434898 417846 435134
rect 448330 435218 448566 435454
rect 448330 434898 448566 435134
rect 479050 435218 479286 435454
rect 479050 434898 479286 435134
rect 509770 435218 510006 435454
rect 509770 434898 510006 435134
rect 540490 435218 540726 435454
rect 540490 434898 540726 435134
rect 33610 417218 33846 417454
rect 33610 416898 33846 417134
rect 64330 417218 64566 417454
rect 64330 416898 64566 417134
rect 95050 417218 95286 417454
rect 95050 416898 95286 417134
rect 125770 417218 126006 417454
rect 125770 416898 126006 417134
rect 156490 417218 156726 417454
rect 156490 416898 156726 417134
rect 187210 417218 187446 417454
rect 187210 416898 187446 417134
rect 217930 417218 218166 417454
rect 217930 416898 218166 417134
rect 248650 417218 248886 417454
rect 248650 416898 248886 417134
rect 279370 417218 279606 417454
rect 279370 416898 279606 417134
rect 310090 417218 310326 417454
rect 310090 416898 310326 417134
rect 340810 417218 341046 417454
rect 340810 416898 341046 417134
rect 371530 417218 371766 417454
rect 371530 416898 371766 417134
rect 402250 417218 402486 417454
rect 402250 416898 402486 417134
rect 432970 417218 433206 417454
rect 432970 416898 433206 417134
rect 463690 417218 463926 417454
rect 463690 416898 463926 417134
rect 494410 417218 494646 417454
rect 494410 416898 494646 417134
rect 525130 417218 525366 417454
rect 525130 416898 525366 417134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 18250 399218 18486 399454
rect 18250 398898 18486 399134
rect 48970 399218 49206 399454
rect 48970 398898 49206 399134
rect 79690 399218 79926 399454
rect 79690 398898 79926 399134
rect 110410 399218 110646 399454
rect 110410 398898 110646 399134
rect 141130 399218 141366 399454
rect 141130 398898 141366 399134
rect 171850 399218 172086 399454
rect 171850 398898 172086 399134
rect 202570 399218 202806 399454
rect 202570 398898 202806 399134
rect 233290 399218 233526 399454
rect 233290 398898 233526 399134
rect 264010 399218 264246 399454
rect 264010 398898 264246 399134
rect 294730 399218 294966 399454
rect 294730 398898 294966 399134
rect 325450 399218 325686 399454
rect 325450 398898 325686 399134
rect 356170 399218 356406 399454
rect 356170 398898 356406 399134
rect 386890 399218 387126 399454
rect 386890 398898 387126 399134
rect 417610 399218 417846 399454
rect 417610 398898 417846 399134
rect 448330 399218 448566 399454
rect 448330 398898 448566 399134
rect 479050 399218 479286 399454
rect 479050 398898 479286 399134
rect 509770 399218 510006 399454
rect 509770 398898 510006 399134
rect 540490 399218 540726 399454
rect 540490 398898 540726 399134
rect 33610 381218 33846 381454
rect 33610 380898 33846 381134
rect 64330 381218 64566 381454
rect 64330 380898 64566 381134
rect 95050 381218 95286 381454
rect 95050 380898 95286 381134
rect 125770 381218 126006 381454
rect 125770 380898 126006 381134
rect 156490 381218 156726 381454
rect 156490 380898 156726 381134
rect 187210 381218 187446 381454
rect 187210 380898 187446 381134
rect 217930 381218 218166 381454
rect 217930 380898 218166 381134
rect 248650 381218 248886 381454
rect 248650 380898 248886 381134
rect 279370 381218 279606 381454
rect 279370 380898 279606 381134
rect 310090 381218 310326 381454
rect 310090 380898 310326 381134
rect 340810 381218 341046 381454
rect 340810 380898 341046 381134
rect 371530 381218 371766 381454
rect 371530 380898 371766 381134
rect 402250 381218 402486 381454
rect 402250 380898 402486 381134
rect 432970 381218 433206 381454
rect 432970 380898 433206 381134
rect 463690 381218 463926 381454
rect 463690 380898 463926 381134
rect 494410 381218 494646 381454
rect 494410 380898 494646 381134
rect 525130 381218 525366 381454
rect 525130 380898 525366 381134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 18250 363218 18486 363454
rect 18250 362898 18486 363134
rect 48970 363218 49206 363454
rect 48970 362898 49206 363134
rect 79690 363218 79926 363454
rect 79690 362898 79926 363134
rect 110410 363218 110646 363454
rect 110410 362898 110646 363134
rect 141130 363218 141366 363454
rect 141130 362898 141366 363134
rect 171850 363218 172086 363454
rect 171850 362898 172086 363134
rect 202570 363218 202806 363454
rect 202570 362898 202806 363134
rect 233290 363218 233526 363454
rect 233290 362898 233526 363134
rect 264010 363218 264246 363454
rect 264010 362898 264246 363134
rect 294730 363218 294966 363454
rect 294730 362898 294966 363134
rect 325450 363218 325686 363454
rect 325450 362898 325686 363134
rect 356170 363218 356406 363454
rect 356170 362898 356406 363134
rect 386890 363218 387126 363454
rect 386890 362898 387126 363134
rect 417610 363218 417846 363454
rect 417610 362898 417846 363134
rect 448330 363218 448566 363454
rect 448330 362898 448566 363134
rect 479050 363218 479286 363454
rect 479050 362898 479286 363134
rect 509770 363218 510006 363454
rect 509770 362898 510006 363134
rect 540490 363218 540726 363454
rect 540490 362898 540726 363134
rect 33610 345218 33846 345454
rect 33610 344898 33846 345134
rect 64330 345218 64566 345454
rect 64330 344898 64566 345134
rect 95050 345218 95286 345454
rect 95050 344898 95286 345134
rect 125770 345218 126006 345454
rect 125770 344898 126006 345134
rect 156490 345218 156726 345454
rect 156490 344898 156726 345134
rect 187210 345218 187446 345454
rect 187210 344898 187446 345134
rect 217930 345218 218166 345454
rect 217930 344898 218166 345134
rect 248650 345218 248886 345454
rect 248650 344898 248886 345134
rect 279370 345218 279606 345454
rect 279370 344898 279606 345134
rect 310090 345218 310326 345454
rect 310090 344898 310326 345134
rect 340810 345218 341046 345454
rect 340810 344898 341046 345134
rect 371530 345218 371766 345454
rect 371530 344898 371766 345134
rect 402250 345218 402486 345454
rect 402250 344898 402486 345134
rect 432970 345218 433206 345454
rect 432970 344898 433206 345134
rect 463690 345218 463926 345454
rect 463690 344898 463926 345134
rect 494410 345218 494646 345454
rect 494410 344898 494646 345134
rect 525130 345218 525366 345454
rect 525130 344898 525366 345134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 18250 327218 18486 327454
rect 18250 326898 18486 327134
rect 48970 327218 49206 327454
rect 48970 326898 49206 327134
rect 79690 327218 79926 327454
rect 79690 326898 79926 327134
rect 110410 327218 110646 327454
rect 110410 326898 110646 327134
rect 141130 327218 141366 327454
rect 141130 326898 141366 327134
rect 171850 327218 172086 327454
rect 171850 326898 172086 327134
rect 202570 327218 202806 327454
rect 202570 326898 202806 327134
rect 233290 327218 233526 327454
rect 233290 326898 233526 327134
rect 264010 327218 264246 327454
rect 264010 326898 264246 327134
rect 294730 327218 294966 327454
rect 294730 326898 294966 327134
rect 325450 327218 325686 327454
rect 325450 326898 325686 327134
rect 356170 327218 356406 327454
rect 356170 326898 356406 327134
rect 386890 327218 387126 327454
rect 386890 326898 387126 327134
rect 417610 327218 417846 327454
rect 417610 326898 417846 327134
rect 448330 327218 448566 327454
rect 448330 326898 448566 327134
rect 479050 327218 479286 327454
rect 479050 326898 479286 327134
rect 509770 327218 510006 327454
rect 509770 326898 510006 327134
rect 540490 327218 540726 327454
rect 540490 326898 540726 327134
rect 33610 309218 33846 309454
rect 33610 308898 33846 309134
rect 64330 309218 64566 309454
rect 64330 308898 64566 309134
rect 95050 309218 95286 309454
rect 95050 308898 95286 309134
rect 125770 309218 126006 309454
rect 125770 308898 126006 309134
rect 156490 309218 156726 309454
rect 156490 308898 156726 309134
rect 187210 309218 187446 309454
rect 187210 308898 187446 309134
rect 217930 309218 218166 309454
rect 217930 308898 218166 309134
rect 248650 309218 248886 309454
rect 248650 308898 248886 309134
rect 279370 309218 279606 309454
rect 279370 308898 279606 309134
rect 310090 309218 310326 309454
rect 310090 308898 310326 309134
rect 340810 309218 341046 309454
rect 340810 308898 341046 309134
rect 371530 309218 371766 309454
rect 371530 308898 371766 309134
rect 402250 309218 402486 309454
rect 402250 308898 402486 309134
rect 432970 309218 433206 309454
rect 432970 308898 433206 309134
rect 463690 309218 463926 309454
rect 463690 308898 463926 309134
rect 494410 309218 494646 309454
rect 494410 308898 494646 309134
rect 525130 309218 525366 309454
rect 525130 308898 525366 309134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 18250 291218 18486 291454
rect 18250 290898 18486 291134
rect 48970 291218 49206 291454
rect 48970 290898 49206 291134
rect 79690 291218 79926 291454
rect 79690 290898 79926 291134
rect 110410 291218 110646 291454
rect 110410 290898 110646 291134
rect 141130 291218 141366 291454
rect 141130 290898 141366 291134
rect 171850 291218 172086 291454
rect 171850 290898 172086 291134
rect 202570 291218 202806 291454
rect 202570 290898 202806 291134
rect 233290 291218 233526 291454
rect 233290 290898 233526 291134
rect 264010 291218 264246 291454
rect 264010 290898 264246 291134
rect 294730 291218 294966 291454
rect 294730 290898 294966 291134
rect 325450 291218 325686 291454
rect 325450 290898 325686 291134
rect 356170 291218 356406 291454
rect 356170 290898 356406 291134
rect 386890 291218 387126 291454
rect 386890 290898 387126 291134
rect 417610 291218 417846 291454
rect 417610 290898 417846 291134
rect 448330 291218 448566 291454
rect 448330 290898 448566 291134
rect 479050 291218 479286 291454
rect 479050 290898 479286 291134
rect 509770 291218 510006 291454
rect 509770 290898 510006 291134
rect 540490 291218 540726 291454
rect 540490 290898 540726 291134
rect 33610 273218 33846 273454
rect 33610 272898 33846 273134
rect 64330 273218 64566 273454
rect 64330 272898 64566 273134
rect 95050 273218 95286 273454
rect 95050 272898 95286 273134
rect 125770 273218 126006 273454
rect 125770 272898 126006 273134
rect 156490 273218 156726 273454
rect 156490 272898 156726 273134
rect 187210 273218 187446 273454
rect 187210 272898 187446 273134
rect 217930 273218 218166 273454
rect 217930 272898 218166 273134
rect 248650 273218 248886 273454
rect 248650 272898 248886 273134
rect 279370 273218 279606 273454
rect 279370 272898 279606 273134
rect 310090 273218 310326 273454
rect 310090 272898 310326 273134
rect 340810 273218 341046 273454
rect 340810 272898 341046 273134
rect 371530 273218 371766 273454
rect 371530 272898 371766 273134
rect 402250 273218 402486 273454
rect 402250 272898 402486 273134
rect 432970 273218 433206 273454
rect 432970 272898 433206 273134
rect 463690 273218 463926 273454
rect 463690 272898 463926 273134
rect 494410 273218 494646 273454
rect 494410 272898 494646 273134
rect 525130 273218 525366 273454
rect 525130 272898 525366 273134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 18250 255218 18486 255454
rect 18250 254898 18486 255134
rect 48970 255218 49206 255454
rect 48970 254898 49206 255134
rect 79690 255218 79926 255454
rect 79690 254898 79926 255134
rect 110410 255218 110646 255454
rect 110410 254898 110646 255134
rect 141130 255218 141366 255454
rect 141130 254898 141366 255134
rect 171850 255218 172086 255454
rect 171850 254898 172086 255134
rect 202570 255218 202806 255454
rect 202570 254898 202806 255134
rect 233290 255218 233526 255454
rect 233290 254898 233526 255134
rect 264010 255218 264246 255454
rect 264010 254898 264246 255134
rect 294730 255218 294966 255454
rect 294730 254898 294966 255134
rect 325450 255218 325686 255454
rect 325450 254898 325686 255134
rect 356170 255218 356406 255454
rect 356170 254898 356406 255134
rect 386890 255218 387126 255454
rect 386890 254898 387126 255134
rect 417610 255218 417846 255454
rect 417610 254898 417846 255134
rect 448330 255218 448566 255454
rect 448330 254898 448566 255134
rect 479050 255218 479286 255454
rect 479050 254898 479286 255134
rect 509770 255218 510006 255454
rect 509770 254898 510006 255134
rect 540490 255218 540726 255454
rect 540490 254898 540726 255134
rect 33610 237218 33846 237454
rect 33610 236898 33846 237134
rect 64330 237218 64566 237454
rect 64330 236898 64566 237134
rect 95050 237218 95286 237454
rect 95050 236898 95286 237134
rect 125770 237218 126006 237454
rect 125770 236898 126006 237134
rect 156490 237218 156726 237454
rect 156490 236898 156726 237134
rect 187210 237218 187446 237454
rect 187210 236898 187446 237134
rect 217930 237218 218166 237454
rect 217930 236898 218166 237134
rect 248650 237218 248886 237454
rect 248650 236898 248886 237134
rect 279370 237218 279606 237454
rect 279370 236898 279606 237134
rect 310090 237218 310326 237454
rect 310090 236898 310326 237134
rect 340810 237218 341046 237454
rect 340810 236898 341046 237134
rect 371530 237218 371766 237454
rect 371530 236898 371766 237134
rect 402250 237218 402486 237454
rect 402250 236898 402486 237134
rect 432970 237218 433206 237454
rect 432970 236898 433206 237134
rect 463690 237218 463926 237454
rect 463690 236898 463926 237134
rect 494410 237218 494646 237454
rect 494410 236898 494646 237134
rect 525130 237218 525366 237454
rect 525130 236898 525366 237134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 18250 219218 18486 219454
rect 18250 218898 18486 219134
rect 48970 219218 49206 219454
rect 48970 218898 49206 219134
rect 79690 219218 79926 219454
rect 79690 218898 79926 219134
rect 110410 219218 110646 219454
rect 110410 218898 110646 219134
rect 141130 219218 141366 219454
rect 141130 218898 141366 219134
rect 171850 219218 172086 219454
rect 171850 218898 172086 219134
rect 202570 219218 202806 219454
rect 202570 218898 202806 219134
rect 233290 219218 233526 219454
rect 233290 218898 233526 219134
rect 264010 219218 264246 219454
rect 264010 218898 264246 219134
rect 294730 219218 294966 219454
rect 294730 218898 294966 219134
rect 325450 219218 325686 219454
rect 325450 218898 325686 219134
rect 356170 219218 356406 219454
rect 356170 218898 356406 219134
rect 386890 219218 387126 219454
rect 386890 218898 387126 219134
rect 417610 219218 417846 219454
rect 417610 218898 417846 219134
rect 448330 219218 448566 219454
rect 448330 218898 448566 219134
rect 479050 219218 479286 219454
rect 479050 218898 479286 219134
rect 509770 219218 510006 219454
rect 509770 218898 510006 219134
rect 540490 219218 540726 219454
rect 540490 218898 540726 219134
rect 33610 201218 33846 201454
rect 33610 200898 33846 201134
rect 64330 201218 64566 201454
rect 64330 200898 64566 201134
rect 95050 201218 95286 201454
rect 95050 200898 95286 201134
rect 125770 201218 126006 201454
rect 125770 200898 126006 201134
rect 156490 201218 156726 201454
rect 156490 200898 156726 201134
rect 187210 201218 187446 201454
rect 187210 200898 187446 201134
rect 217930 201218 218166 201454
rect 217930 200898 218166 201134
rect 248650 201218 248886 201454
rect 248650 200898 248886 201134
rect 279370 201218 279606 201454
rect 279370 200898 279606 201134
rect 310090 201218 310326 201454
rect 310090 200898 310326 201134
rect 340810 201218 341046 201454
rect 340810 200898 341046 201134
rect 371530 201218 371766 201454
rect 371530 200898 371766 201134
rect 402250 201218 402486 201454
rect 402250 200898 402486 201134
rect 432970 201218 433206 201454
rect 432970 200898 433206 201134
rect 463690 201218 463926 201454
rect 463690 200898 463926 201134
rect 494410 201218 494646 201454
rect 494410 200898 494646 201134
rect 525130 201218 525366 201454
rect 525130 200898 525366 201134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 18250 183218 18486 183454
rect 18250 182898 18486 183134
rect 48970 183218 49206 183454
rect 48970 182898 49206 183134
rect 79690 183218 79926 183454
rect 79690 182898 79926 183134
rect 110410 183218 110646 183454
rect 110410 182898 110646 183134
rect 141130 183218 141366 183454
rect 141130 182898 141366 183134
rect 171850 183218 172086 183454
rect 171850 182898 172086 183134
rect 202570 183218 202806 183454
rect 202570 182898 202806 183134
rect 233290 183218 233526 183454
rect 233290 182898 233526 183134
rect 264010 183218 264246 183454
rect 264010 182898 264246 183134
rect 294730 183218 294966 183454
rect 294730 182898 294966 183134
rect 325450 183218 325686 183454
rect 325450 182898 325686 183134
rect 356170 183218 356406 183454
rect 356170 182898 356406 183134
rect 386890 183218 387126 183454
rect 386890 182898 387126 183134
rect 417610 183218 417846 183454
rect 417610 182898 417846 183134
rect 448330 183218 448566 183454
rect 448330 182898 448566 183134
rect 479050 183218 479286 183454
rect 479050 182898 479286 183134
rect 509770 183218 510006 183454
rect 509770 182898 510006 183134
rect 540490 183218 540726 183454
rect 540490 182898 540726 183134
rect 33610 165218 33846 165454
rect 33610 164898 33846 165134
rect 64330 165218 64566 165454
rect 64330 164898 64566 165134
rect 95050 165218 95286 165454
rect 95050 164898 95286 165134
rect 125770 165218 126006 165454
rect 125770 164898 126006 165134
rect 156490 165218 156726 165454
rect 156490 164898 156726 165134
rect 187210 165218 187446 165454
rect 187210 164898 187446 165134
rect 217930 165218 218166 165454
rect 217930 164898 218166 165134
rect 248650 165218 248886 165454
rect 248650 164898 248886 165134
rect 279370 165218 279606 165454
rect 279370 164898 279606 165134
rect 310090 165218 310326 165454
rect 310090 164898 310326 165134
rect 340810 165218 341046 165454
rect 340810 164898 341046 165134
rect 371530 165218 371766 165454
rect 371530 164898 371766 165134
rect 402250 165218 402486 165454
rect 402250 164898 402486 165134
rect 432970 165218 433206 165454
rect 432970 164898 433206 165134
rect 463690 165218 463926 165454
rect 463690 164898 463926 165134
rect 494410 165218 494646 165454
rect 494410 164898 494646 165134
rect 525130 165218 525366 165454
rect 525130 164898 525366 165134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 18250 147218 18486 147454
rect 18250 146898 18486 147134
rect 48970 147218 49206 147454
rect 48970 146898 49206 147134
rect 79690 147218 79926 147454
rect 79690 146898 79926 147134
rect 110410 147218 110646 147454
rect 110410 146898 110646 147134
rect 141130 147218 141366 147454
rect 141130 146898 141366 147134
rect 171850 147218 172086 147454
rect 171850 146898 172086 147134
rect 202570 147218 202806 147454
rect 202570 146898 202806 147134
rect 233290 147218 233526 147454
rect 233290 146898 233526 147134
rect 264010 147218 264246 147454
rect 264010 146898 264246 147134
rect 294730 147218 294966 147454
rect 294730 146898 294966 147134
rect 325450 147218 325686 147454
rect 325450 146898 325686 147134
rect 356170 147218 356406 147454
rect 356170 146898 356406 147134
rect 386890 147218 387126 147454
rect 386890 146898 387126 147134
rect 417610 147218 417846 147454
rect 417610 146898 417846 147134
rect 448330 147218 448566 147454
rect 448330 146898 448566 147134
rect 479050 147218 479286 147454
rect 479050 146898 479286 147134
rect 509770 147218 510006 147454
rect 509770 146898 510006 147134
rect 540490 147218 540726 147454
rect 540490 146898 540726 147134
rect 33610 129218 33846 129454
rect 33610 128898 33846 129134
rect 64330 129218 64566 129454
rect 64330 128898 64566 129134
rect 95050 129218 95286 129454
rect 95050 128898 95286 129134
rect 125770 129218 126006 129454
rect 125770 128898 126006 129134
rect 156490 129218 156726 129454
rect 156490 128898 156726 129134
rect 187210 129218 187446 129454
rect 187210 128898 187446 129134
rect 217930 129218 218166 129454
rect 217930 128898 218166 129134
rect 248650 129218 248886 129454
rect 248650 128898 248886 129134
rect 279370 129218 279606 129454
rect 279370 128898 279606 129134
rect 310090 129218 310326 129454
rect 310090 128898 310326 129134
rect 340810 129218 341046 129454
rect 340810 128898 341046 129134
rect 371530 129218 371766 129454
rect 371530 128898 371766 129134
rect 402250 129218 402486 129454
rect 402250 128898 402486 129134
rect 432970 129218 433206 129454
rect 432970 128898 433206 129134
rect 463690 129218 463926 129454
rect 463690 128898 463926 129134
rect 494410 129218 494646 129454
rect 494410 128898 494646 129134
rect 525130 129218 525366 129454
rect 525130 128898 525366 129134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 18250 111218 18486 111454
rect 18250 110898 18486 111134
rect 48970 111218 49206 111454
rect 48970 110898 49206 111134
rect 79690 111218 79926 111454
rect 79690 110898 79926 111134
rect 110410 111218 110646 111454
rect 110410 110898 110646 111134
rect 141130 111218 141366 111454
rect 141130 110898 141366 111134
rect 171850 111218 172086 111454
rect 171850 110898 172086 111134
rect 202570 111218 202806 111454
rect 202570 110898 202806 111134
rect 233290 111218 233526 111454
rect 233290 110898 233526 111134
rect 264010 111218 264246 111454
rect 264010 110898 264246 111134
rect 294730 111218 294966 111454
rect 294730 110898 294966 111134
rect 325450 111218 325686 111454
rect 325450 110898 325686 111134
rect 356170 111218 356406 111454
rect 356170 110898 356406 111134
rect 386890 111218 387126 111454
rect 386890 110898 387126 111134
rect 417610 111218 417846 111454
rect 417610 110898 417846 111134
rect 448330 111218 448566 111454
rect 448330 110898 448566 111134
rect 479050 111218 479286 111454
rect 479050 110898 479286 111134
rect 509770 111218 510006 111454
rect 509770 110898 510006 111134
rect 540490 111218 540726 111454
rect 540490 110898 540726 111134
rect 33610 93218 33846 93454
rect 33610 92898 33846 93134
rect 64330 93218 64566 93454
rect 64330 92898 64566 93134
rect 95050 93218 95286 93454
rect 95050 92898 95286 93134
rect 125770 93218 126006 93454
rect 125770 92898 126006 93134
rect 156490 93218 156726 93454
rect 156490 92898 156726 93134
rect 187210 93218 187446 93454
rect 187210 92898 187446 93134
rect 217930 93218 218166 93454
rect 217930 92898 218166 93134
rect 248650 93218 248886 93454
rect 248650 92898 248886 93134
rect 279370 93218 279606 93454
rect 279370 92898 279606 93134
rect 310090 93218 310326 93454
rect 310090 92898 310326 93134
rect 340810 93218 341046 93454
rect 340810 92898 341046 93134
rect 371530 93218 371766 93454
rect 371530 92898 371766 93134
rect 402250 93218 402486 93454
rect 402250 92898 402486 93134
rect 432970 93218 433206 93454
rect 432970 92898 433206 93134
rect 463690 93218 463926 93454
rect 463690 92898 463926 93134
rect 494410 93218 494646 93454
rect 494410 92898 494646 93134
rect 525130 93218 525366 93454
rect 525130 92898 525366 93134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 18250 75218 18486 75454
rect 18250 74898 18486 75134
rect 48970 75218 49206 75454
rect 48970 74898 49206 75134
rect 79690 75218 79926 75454
rect 79690 74898 79926 75134
rect 110410 75218 110646 75454
rect 110410 74898 110646 75134
rect 141130 75218 141366 75454
rect 141130 74898 141366 75134
rect 171850 75218 172086 75454
rect 171850 74898 172086 75134
rect 202570 75218 202806 75454
rect 202570 74898 202806 75134
rect 233290 75218 233526 75454
rect 233290 74898 233526 75134
rect 264010 75218 264246 75454
rect 264010 74898 264246 75134
rect 294730 75218 294966 75454
rect 294730 74898 294966 75134
rect 325450 75218 325686 75454
rect 325450 74898 325686 75134
rect 356170 75218 356406 75454
rect 356170 74898 356406 75134
rect 386890 75218 387126 75454
rect 386890 74898 387126 75134
rect 417610 75218 417846 75454
rect 417610 74898 417846 75134
rect 448330 75218 448566 75454
rect 448330 74898 448566 75134
rect 479050 75218 479286 75454
rect 479050 74898 479286 75134
rect 509770 75218 510006 75454
rect 509770 74898 510006 75134
rect 540490 75218 540726 75454
rect 540490 74898 540726 75134
rect 33610 57218 33846 57454
rect 33610 56898 33846 57134
rect 64330 57218 64566 57454
rect 64330 56898 64566 57134
rect 95050 57218 95286 57454
rect 95050 56898 95286 57134
rect 125770 57218 126006 57454
rect 125770 56898 126006 57134
rect 156490 57218 156726 57454
rect 156490 56898 156726 57134
rect 187210 57218 187446 57454
rect 187210 56898 187446 57134
rect 217930 57218 218166 57454
rect 217930 56898 218166 57134
rect 248650 57218 248886 57454
rect 248650 56898 248886 57134
rect 279370 57218 279606 57454
rect 279370 56898 279606 57134
rect 310090 57218 310326 57454
rect 310090 56898 310326 57134
rect 340810 57218 341046 57454
rect 340810 56898 341046 57134
rect 371530 57218 371766 57454
rect 371530 56898 371766 57134
rect 402250 57218 402486 57454
rect 402250 56898 402486 57134
rect 432970 57218 433206 57454
rect 432970 56898 433206 57134
rect 463690 57218 463926 57454
rect 463690 56898 463926 57134
rect 494410 57218 494646 57454
rect 494410 56898 494646 57134
rect 525130 57218 525366 57454
rect 525130 56898 525366 57134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 18250 651454
rect 18486 651218 48970 651454
rect 49206 651218 79690 651454
rect 79926 651218 110410 651454
rect 110646 651218 141130 651454
rect 141366 651218 171850 651454
rect 172086 651218 202570 651454
rect 202806 651218 233290 651454
rect 233526 651218 264010 651454
rect 264246 651218 294730 651454
rect 294966 651218 325450 651454
rect 325686 651218 356170 651454
rect 356406 651218 386890 651454
rect 387126 651218 417610 651454
rect 417846 651218 448330 651454
rect 448566 651218 479050 651454
rect 479286 651218 509770 651454
rect 510006 651218 540490 651454
rect 540726 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 18250 651134
rect 18486 650898 48970 651134
rect 49206 650898 79690 651134
rect 79926 650898 110410 651134
rect 110646 650898 141130 651134
rect 141366 650898 171850 651134
rect 172086 650898 202570 651134
rect 202806 650898 233290 651134
rect 233526 650898 264010 651134
rect 264246 650898 294730 651134
rect 294966 650898 325450 651134
rect 325686 650898 356170 651134
rect 356406 650898 386890 651134
rect 387126 650898 417610 651134
rect 417846 650898 448330 651134
rect 448566 650898 479050 651134
rect 479286 650898 509770 651134
rect 510006 650898 540490 651134
rect 540726 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 33610 633454
rect 33846 633218 64330 633454
rect 64566 633218 95050 633454
rect 95286 633218 125770 633454
rect 126006 633218 156490 633454
rect 156726 633218 187210 633454
rect 187446 633218 217930 633454
rect 218166 633218 248650 633454
rect 248886 633218 279370 633454
rect 279606 633218 310090 633454
rect 310326 633218 340810 633454
rect 341046 633218 371530 633454
rect 371766 633218 402250 633454
rect 402486 633218 432970 633454
rect 433206 633218 463690 633454
rect 463926 633218 494410 633454
rect 494646 633218 525130 633454
rect 525366 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 33610 633134
rect 33846 632898 64330 633134
rect 64566 632898 95050 633134
rect 95286 632898 125770 633134
rect 126006 632898 156490 633134
rect 156726 632898 187210 633134
rect 187446 632898 217930 633134
rect 218166 632898 248650 633134
rect 248886 632898 279370 633134
rect 279606 632898 310090 633134
rect 310326 632898 340810 633134
rect 341046 632898 371530 633134
rect 371766 632898 402250 633134
rect 402486 632898 432970 633134
rect 433206 632898 463690 633134
rect 463926 632898 494410 633134
rect 494646 632898 525130 633134
rect 525366 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 18250 615454
rect 18486 615218 48970 615454
rect 49206 615218 79690 615454
rect 79926 615218 110410 615454
rect 110646 615218 141130 615454
rect 141366 615218 171850 615454
rect 172086 615218 202570 615454
rect 202806 615218 233290 615454
rect 233526 615218 264010 615454
rect 264246 615218 294730 615454
rect 294966 615218 325450 615454
rect 325686 615218 356170 615454
rect 356406 615218 386890 615454
rect 387126 615218 417610 615454
rect 417846 615218 448330 615454
rect 448566 615218 479050 615454
rect 479286 615218 509770 615454
rect 510006 615218 540490 615454
rect 540726 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 18250 615134
rect 18486 614898 48970 615134
rect 49206 614898 79690 615134
rect 79926 614898 110410 615134
rect 110646 614898 141130 615134
rect 141366 614898 171850 615134
rect 172086 614898 202570 615134
rect 202806 614898 233290 615134
rect 233526 614898 264010 615134
rect 264246 614898 294730 615134
rect 294966 614898 325450 615134
rect 325686 614898 356170 615134
rect 356406 614898 386890 615134
rect 387126 614898 417610 615134
rect 417846 614898 448330 615134
rect 448566 614898 479050 615134
rect 479286 614898 509770 615134
rect 510006 614898 540490 615134
rect 540726 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 33610 597454
rect 33846 597218 64330 597454
rect 64566 597218 95050 597454
rect 95286 597218 125770 597454
rect 126006 597218 156490 597454
rect 156726 597218 187210 597454
rect 187446 597218 217930 597454
rect 218166 597218 248650 597454
rect 248886 597218 279370 597454
rect 279606 597218 310090 597454
rect 310326 597218 340810 597454
rect 341046 597218 371530 597454
rect 371766 597218 402250 597454
rect 402486 597218 432970 597454
rect 433206 597218 463690 597454
rect 463926 597218 494410 597454
rect 494646 597218 525130 597454
rect 525366 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 33610 597134
rect 33846 596898 64330 597134
rect 64566 596898 95050 597134
rect 95286 596898 125770 597134
rect 126006 596898 156490 597134
rect 156726 596898 187210 597134
rect 187446 596898 217930 597134
rect 218166 596898 248650 597134
rect 248886 596898 279370 597134
rect 279606 596898 310090 597134
rect 310326 596898 340810 597134
rect 341046 596898 371530 597134
rect 371766 596898 402250 597134
rect 402486 596898 432970 597134
rect 433206 596898 463690 597134
rect 463926 596898 494410 597134
rect 494646 596898 525130 597134
rect 525366 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 18250 579454
rect 18486 579218 48970 579454
rect 49206 579218 79690 579454
rect 79926 579218 110410 579454
rect 110646 579218 141130 579454
rect 141366 579218 171850 579454
rect 172086 579218 202570 579454
rect 202806 579218 233290 579454
rect 233526 579218 264010 579454
rect 264246 579218 294730 579454
rect 294966 579218 325450 579454
rect 325686 579218 356170 579454
rect 356406 579218 386890 579454
rect 387126 579218 417610 579454
rect 417846 579218 448330 579454
rect 448566 579218 479050 579454
rect 479286 579218 509770 579454
rect 510006 579218 540490 579454
rect 540726 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 18250 579134
rect 18486 578898 48970 579134
rect 49206 578898 79690 579134
rect 79926 578898 110410 579134
rect 110646 578898 141130 579134
rect 141366 578898 171850 579134
rect 172086 578898 202570 579134
rect 202806 578898 233290 579134
rect 233526 578898 264010 579134
rect 264246 578898 294730 579134
rect 294966 578898 325450 579134
rect 325686 578898 356170 579134
rect 356406 578898 386890 579134
rect 387126 578898 417610 579134
rect 417846 578898 448330 579134
rect 448566 578898 479050 579134
rect 479286 578898 509770 579134
rect 510006 578898 540490 579134
rect 540726 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 33610 561454
rect 33846 561218 64330 561454
rect 64566 561218 95050 561454
rect 95286 561218 125770 561454
rect 126006 561218 156490 561454
rect 156726 561218 187210 561454
rect 187446 561218 217930 561454
rect 218166 561218 248650 561454
rect 248886 561218 279370 561454
rect 279606 561218 310090 561454
rect 310326 561218 340810 561454
rect 341046 561218 371530 561454
rect 371766 561218 402250 561454
rect 402486 561218 432970 561454
rect 433206 561218 463690 561454
rect 463926 561218 494410 561454
rect 494646 561218 525130 561454
rect 525366 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 33610 561134
rect 33846 560898 64330 561134
rect 64566 560898 95050 561134
rect 95286 560898 125770 561134
rect 126006 560898 156490 561134
rect 156726 560898 187210 561134
rect 187446 560898 217930 561134
rect 218166 560898 248650 561134
rect 248886 560898 279370 561134
rect 279606 560898 310090 561134
rect 310326 560898 340810 561134
rect 341046 560898 371530 561134
rect 371766 560898 402250 561134
rect 402486 560898 432970 561134
rect 433206 560898 463690 561134
rect 463926 560898 494410 561134
rect 494646 560898 525130 561134
rect 525366 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 18250 543454
rect 18486 543218 48970 543454
rect 49206 543218 79690 543454
rect 79926 543218 110410 543454
rect 110646 543218 141130 543454
rect 141366 543218 171850 543454
rect 172086 543218 202570 543454
rect 202806 543218 233290 543454
rect 233526 543218 264010 543454
rect 264246 543218 294730 543454
rect 294966 543218 325450 543454
rect 325686 543218 356170 543454
rect 356406 543218 386890 543454
rect 387126 543218 417610 543454
rect 417846 543218 448330 543454
rect 448566 543218 479050 543454
rect 479286 543218 509770 543454
rect 510006 543218 540490 543454
rect 540726 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 18250 543134
rect 18486 542898 48970 543134
rect 49206 542898 79690 543134
rect 79926 542898 110410 543134
rect 110646 542898 141130 543134
rect 141366 542898 171850 543134
rect 172086 542898 202570 543134
rect 202806 542898 233290 543134
rect 233526 542898 264010 543134
rect 264246 542898 294730 543134
rect 294966 542898 325450 543134
rect 325686 542898 356170 543134
rect 356406 542898 386890 543134
rect 387126 542898 417610 543134
rect 417846 542898 448330 543134
rect 448566 542898 479050 543134
rect 479286 542898 509770 543134
rect 510006 542898 540490 543134
rect 540726 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 33610 525454
rect 33846 525218 64330 525454
rect 64566 525218 95050 525454
rect 95286 525218 125770 525454
rect 126006 525218 156490 525454
rect 156726 525218 187210 525454
rect 187446 525218 217930 525454
rect 218166 525218 248650 525454
rect 248886 525218 279370 525454
rect 279606 525218 310090 525454
rect 310326 525218 340810 525454
rect 341046 525218 371530 525454
rect 371766 525218 402250 525454
rect 402486 525218 432970 525454
rect 433206 525218 463690 525454
rect 463926 525218 494410 525454
rect 494646 525218 525130 525454
rect 525366 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 33610 525134
rect 33846 524898 64330 525134
rect 64566 524898 95050 525134
rect 95286 524898 125770 525134
rect 126006 524898 156490 525134
rect 156726 524898 187210 525134
rect 187446 524898 217930 525134
rect 218166 524898 248650 525134
rect 248886 524898 279370 525134
rect 279606 524898 310090 525134
rect 310326 524898 340810 525134
rect 341046 524898 371530 525134
rect 371766 524898 402250 525134
rect 402486 524898 432970 525134
rect 433206 524898 463690 525134
rect 463926 524898 494410 525134
rect 494646 524898 525130 525134
rect 525366 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 18250 507454
rect 18486 507218 48970 507454
rect 49206 507218 79690 507454
rect 79926 507218 110410 507454
rect 110646 507218 141130 507454
rect 141366 507218 171850 507454
rect 172086 507218 202570 507454
rect 202806 507218 233290 507454
rect 233526 507218 264010 507454
rect 264246 507218 294730 507454
rect 294966 507218 325450 507454
rect 325686 507218 356170 507454
rect 356406 507218 386890 507454
rect 387126 507218 417610 507454
rect 417846 507218 448330 507454
rect 448566 507218 479050 507454
rect 479286 507218 509770 507454
rect 510006 507218 540490 507454
rect 540726 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 18250 507134
rect 18486 506898 48970 507134
rect 49206 506898 79690 507134
rect 79926 506898 110410 507134
rect 110646 506898 141130 507134
rect 141366 506898 171850 507134
rect 172086 506898 202570 507134
rect 202806 506898 233290 507134
rect 233526 506898 264010 507134
rect 264246 506898 294730 507134
rect 294966 506898 325450 507134
rect 325686 506898 356170 507134
rect 356406 506898 386890 507134
rect 387126 506898 417610 507134
rect 417846 506898 448330 507134
rect 448566 506898 479050 507134
rect 479286 506898 509770 507134
rect 510006 506898 540490 507134
rect 540726 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 33610 489454
rect 33846 489218 64330 489454
rect 64566 489218 95050 489454
rect 95286 489218 125770 489454
rect 126006 489218 156490 489454
rect 156726 489218 187210 489454
rect 187446 489218 217930 489454
rect 218166 489218 248650 489454
rect 248886 489218 279370 489454
rect 279606 489218 310090 489454
rect 310326 489218 340810 489454
rect 341046 489218 371530 489454
rect 371766 489218 402250 489454
rect 402486 489218 432970 489454
rect 433206 489218 463690 489454
rect 463926 489218 494410 489454
rect 494646 489218 525130 489454
rect 525366 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 33610 489134
rect 33846 488898 64330 489134
rect 64566 488898 95050 489134
rect 95286 488898 125770 489134
rect 126006 488898 156490 489134
rect 156726 488898 187210 489134
rect 187446 488898 217930 489134
rect 218166 488898 248650 489134
rect 248886 488898 279370 489134
rect 279606 488898 310090 489134
rect 310326 488898 340810 489134
rect 341046 488898 371530 489134
rect 371766 488898 402250 489134
rect 402486 488898 432970 489134
rect 433206 488898 463690 489134
rect 463926 488898 494410 489134
rect 494646 488898 525130 489134
rect 525366 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 18250 471454
rect 18486 471218 48970 471454
rect 49206 471218 79690 471454
rect 79926 471218 110410 471454
rect 110646 471218 141130 471454
rect 141366 471218 171850 471454
rect 172086 471218 202570 471454
rect 202806 471218 233290 471454
rect 233526 471218 264010 471454
rect 264246 471218 294730 471454
rect 294966 471218 325450 471454
rect 325686 471218 356170 471454
rect 356406 471218 386890 471454
rect 387126 471218 417610 471454
rect 417846 471218 448330 471454
rect 448566 471218 479050 471454
rect 479286 471218 509770 471454
rect 510006 471218 540490 471454
rect 540726 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 18250 471134
rect 18486 470898 48970 471134
rect 49206 470898 79690 471134
rect 79926 470898 110410 471134
rect 110646 470898 141130 471134
rect 141366 470898 171850 471134
rect 172086 470898 202570 471134
rect 202806 470898 233290 471134
rect 233526 470898 264010 471134
rect 264246 470898 294730 471134
rect 294966 470898 325450 471134
rect 325686 470898 356170 471134
rect 356406 470898 386890 471134
rect 387126 470898 417610 471134
rect 417846 470898 448330 471134
rect 448566 470898 479050 471134
rect 479286 470898 509770 471134
rect 510006 470898 540490 471134
rect 540726 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 33610 453454
rect 33846 453218 64330 453454
rect 64566 453218 95050 453454
rect 95286 453218 125770 453454
rect 126006 453218 156490 453454
rect 156726 453218 187210 453454
rect 187446 453218 217930 453454
rect 218166 453218 248650 453454
rect 248886 453218 279370 453454
rect 279606 453218 310090 453454
rect 310326 453218 340810 453454
rect 341046 453218 371530 453454
rect 371766 453218 402250 453454
rect 402486 453218 432970 453454
rect 433206 453218 463690 453454
rect 463926 453218 494410 453454
rect 494646 453218 525130 453454
rect 525366 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 33610 453134
rect 33846 452898 64330 453134
rect 64566 452898 95050 453134
rect 95286 452898 125770 453134
rect 126006 452898 156490 453134
rect 156726 452898 187210 453134
rect 187446 452898 217930 453134
rect 218166 452898 248650 453134
rect 248886 452898 279370 453134
rect 279606 452898 310090 453134
rect 310326 452898 340810 453134
rect 341046 452898 371530 453134
rect 371766 452898 402250 453134
rect 402486 452898 432970 453134
rect 433206 452898 463690 453134
rect 463926 452898 494410 453134
rect 494646 452898 525130 453134
rect 525366 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 18250 435454
rect 18486 435218 48970 435454
rect 49206 435218 79690 435454
rect 79926 435218 110410 435454
rect 110646 435218 141130 435454
rect 141366 435218 171850 435454
rect 172086 435218 202570 435454
rect 202806 435218 233290 435454
rect 233526 435218 264010 435454
rect 264246 435218 294730 435454
rect 294966 435218 325450 435454
rect 325686 435218 356170 435454
rect 356406 435218 386890 435454
rect 387126 435218 417610 435454
rect 417846 435218 448330 435454
rect 448566 435218 479050 435454
rect 479286 435218 509770 435454
rect 510006 435218 540490 435454
rect 540726 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 18250 435134
rect 18486 434898 48970 435134
rect 49206 434898 79690 435134
rect 79926 434898 110410 435134
rect 110646 434898 141130 435134
rect 141366 434898 171850 435134
rect 172086 434898 202570 435134
rect 202806 434898 233290 435134
rect 233526 434898 264010 435134
rect 264246 434898 294730 435134
rect 294966 434898 325450 435134
rect 325686 434898 356170 435134
rect 356406 434898 386890 435134
rect 387126 434898 417610 435134
rect 417846 434898 448330 435134
rect 448566 434898 479050 435134
rect 479286 434898 509770 435134
rect 510006 434898 540490 435134
rect 540726 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 33610 417454
rect 33846 417218 64330 417454
rect 64566 417218 95050 417454
rect 95286 417218 125770 417454
rect 126006 417218 156490 417454
rect 156726 417218 187210 417454
rect 187446 417218 217930 417454
rect 218166 417218 248650 417454
rect 248886 417218 279370 417454
rect 279606 417218 310090 417454
rect 310326 417218 340810 417454
rect 341046 417218 371530 417454
rect 371766 417218 402250 417454
rect 402486 417218 432970 417454
rect 433206 417218 463690 417454
rect 463926 417218 494410 417454
rect 494646 417218 525130 417454
rect 525366 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 33610 417134
rect 33846 416898 64330 417134
rect 64566 416898 95050 417134
rect 95286 416898 125770 417134
rect 126006 416898 156490 417134
rect 156726 416898 187210 417134
rect 187446 416898 217930 417134
rect 218166 416898 248650 417134
rect 248886 416898 279370 417134
rect 279606 416898 310090 417134
rect 310326 416898 340810 417134
rect 341046 416898 371530 417134
rect 371766 416898 402250 417134
rect 402486 416898 432970 417134
rect 433206 416898 463690 417134
rect 463926 416898 494410 417134
rect 494646 416898 525130 417134
rect 525366 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 18250 399454
rect 18486 399218 48970 399454
rect 49206 399218 79690 399454
rect 79926 399218 110410 399454
rect 110646 399218 141130 399454
rect 141366 399218 171850 399454
rect 172086 399218 202570 399454
rect 202806 399218 233290 399454
rect 233526 399218 264010 399454
rect 264246 399218 294730 399454
rect 294966 399218 325450 399454
rect 325686 399218 356170 399454
rect 356406 399218 386890 399454
rect 387126 399218 417610 399454
rect 417846 399218 448330 399454
rect 448566 399218 479050 399454
rect 479286 399218 509770 399454
rect 510006 399218 540490 399454
rect 540726 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 18250 399134
rect 18486 398898 48970 399134
rect 49206 398898 79690 399134
rect 79926 398898 110410 399134
rect 110646 398898 141130 399134
rect 141366 398898 171850 399134
rect 172086 398898 202570 399134
rect 202806 398898 233290 399134
rect 233526 398898 264010 399134
rect 264246 398898 294730 399134
rect 294966 398898 325450 399134
rect 325686 398898 356170 399134
rect 356406 398898 386890 399134
rect 387126 398898 417610 399134
rect 417846 398898 448330 399134
rect 448566 398898 479050 399134
rect 479286 398898 509770 399134
rect 510006 398898 540490 399134
rect 540726 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 33610 381454
rect 33846 381218 64330 381454
rect 64566 381218 95050 381454
rect 95286 381218 125770 381454
rect 126006 381218 156490 381454
rect 156726 381218 187210 381454
rect 187446 381218 217930 381454
rect 218166 381218 248650 381454
rect 248886 381218 279370 381454
rect 279606 381218 310090 381454
rect 310326 381218 340810 381454
rect 341046 381218 371530 381454
rect 371766 381218 402250 381454
rect 402486 381218 432970 381454
rect 433206 381218 463690 381454
rect 463926 381218 494410 381454
rect 494646 381218 525130 381454
rect 525366 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 33610 381134
rect 33846 380898 64330 381134
rect 64566 380898 95050 381134
rect 95286 380898 125770 381134
rect 126006 380898 156490 381134
rect 156726 380898 187210 381134
rect 187446 380898 217930 381134
rect 218166 380898 248650 381134
rect 248886 380898 279370 381134
rect 279606 380898 310090 381134
rect 310326 380898 340810 381134
rect 341046 380898 371530 381134
rect 371766 380898 402250 381134
rect 402486 380898 432970 381134
rect 433206 380898 463690 381134
rect 463926 380898 494410 381134
rect 494646 380898 525130 381134
rect 525366 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 18250 363454
rect 18486 363218 48970 363454
rect 49206 363218 79690 363454
rect 79926 363218 110410 363454
rect 110646 363218 141130 363454
rect 141366 363218 171850 363454
rect 172086 363218 202570 363454
rect 202806 363218 233290 363454
rect 233526 363218 264010 363454
rect 264246 363218 294730 363454
rect 294966 363218 325450 363454
rect 325686 363218 356170 363454
rect 356406 363218 386890 363454
rect 387126 363218 417610 363454
rect 417846 363218 448330 363454
rect 448566 363218 479050 363454
rect 479286 363218 509770 363454
rect 510006 363218 540490 363454
rect 540726 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 18250 363134
rect 18486 362898 48970 363134
rect 49206 362898 79690 363134
rect 79926 362898 110410 363134
rect 110646 362898 141130 363134
rect 141366 362898 171850 363134
rect 172086 362898 202570 363134
rect 202806 362898 233290 363134
rect 233526 362898 264010 363134
rect 264246 362898 294730 363134
rect 294966 362898 325450 363134
rect 325686 362898 356170 363134
rect 356406 362898 386890 363134
rect 387126 362898 417610 363134
rect 417846 362898 448330 363134
rect 448566 362898 479050 363134
rect 479286 362898 509770 363134
rect 510006 362898 540490 363134
rect 540726 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 33610 345454
rect 33846 345218 64330 345454
rect 64566 345218 95050 345454
rect 95286 345218 125770 345454
rect 126006 345218 156490 345454
rect 156726 345218 187210 345454
rect 187446 345218 217930 345454
rect 218166 345218 248650 345454
rect 248886 345218 279370 345454
rect 279606 345218 310090 345454
rect 310326 345218 340810 345454
rect 341046 345218 371530 345454
rect 371766 345218 402250 345454
rect 402486 345218 432970 345454
rect 433206 345218 463690 345454
rect 463926 345218 494410 345454
rect 494646 345218 525130 345454
rect 525366 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 33610 345134
rect 33846 344898 64330 345134
rect 64566 344898 95050 345134
rect 95286 344898 125770 345134
rect 126006 344898 156490 345134
rect 156726 344898 187210 345134
rect 187446 344898 217930 345134
rect 218166 344898 248650 345134
rect 248886 344898 279370 345134
rect 279606 344898 310090 345134
rect 310326 344898 340810 345134
rect 341046 344898 371530 345134
rect 371766 344898 402250 345134
rect 402486 344898 432970 345134
rect 433206 344898 463690 345134
rect 463926 344898 494410 345134
rect 494646 344898 525130 345134
rect 525366 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 18250 327454
rect 18486 327218 48970 327454
rect 49206 327218 79690 327454
rect 79926 327218 110410 327454
rect 110646 327218 141130 327454
rect 141366 327218 171850 327454
rect 172086 327218 202570 327454
rect 202806 327218 233290 327454
rect 233526 327218 264010 327454
rect 264246 327218 294730 327454
rect 294966 327218 325450 327454
rect 325686 327218 356170 327454
rect 356406 327218 386890 327454
rect 387126 327218 417610 327454
rect 417846 327218 448330 327454
rect 448566 327218 479050 327454
rect 479286 327218 509770 327454
rect 510006 327218 540490 327454
rect 540726 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 18250 327134
rect 18486 326898 48970 327134
rect 49206 326898 79690 327134
rect 79926 326898 110410 327134
rect 110646 326898 141130 327134
rect 141366 326898 171850 327134
rect 172086 326898 202570 327134
rect 202806 326898 233290 327134
rect 233526 326898 264010 327134
rect 264246 326898 294730 327134
rect 294966 326898 325450 327134
rect 325686 326898 356170 327134
rect 356406 326898 386890 327134
rect 387126 326898 417610 327134
rect 417846 326898 448330 327134
rect 448566 326898 479050 327134
rect 479286 326898 509770 327134
rect 510006 326898 540490 327134
rect 540726 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 33610 309454
rect 33846 309218 64330 309454
rect 64566 309218 95050 309454
rect 95286 309218 125770 309454
rect 126006 309218 156490 309454
rect 156726 309218 187210 309454
rect 187446 309218 217930 309454
rect 218166 309218 248650 309454
rect 248886 309218 279370 309454
rect 279606 309218 310090 309454
rect 310326 309218 340810 309454
rect 341046 309218 371530 309454
rect 371766 309218 402250 309454
rect 402486 309218 432970 309454
rect 433206 309218 463690 309454
rect 463926 309218 494410 309454
rect 494646 309218 525130 309454
rect 525366 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 33610 309134
rect 33846 308898 64330 309134
rect 64566 308898 95050 309134
rect 95286 308898 125770 309134
rect 126006 308898 156490 309134
rect 156726 308898 187210 309134
rect 187446 308898 217930 309134
rect 218166 308898 248650 309134
rect 248886 308898 279370 309134
rect 279606 308898 310090 309134
rect 310326 308898 340810 309134
rect 341046 308898 371530 309134
rect 371766 308898 402250 309134
rect 402486 308898 432970 309134
rect 433206 308898 463690 309134
rect 463926 308898 494410 309134
rect 494646 308898 525130 309134
rect 525366 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 18250 291454
rect 18486 291218 48970 291454
rect 49206 291218 79690 291454
rect 79926 291218 110410 291454
rect 110646 291218 141130 291454
rect 141366 291218 171850 291454
rect 172086 291218 202570 291454
rect 202806 291218 233290 291454
rect 233526 291218 264010 291454
rect 264246 291218 294730 291454
rect 294966 291218 325450 291454
rect 325686 291218 356170 291454
rect 356406 291218 386890 291454
rect 387126 291218 417610 291454
rect 417846 291218 448330 291454
rect 448566 291218 479050 291454
rect 479286 291218 509770 291454
rect 510006 291218 540490 291454
rect 540726 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 18250 291134
rect 18486 290898 48970 291134
rect 49206 290898 79690 291134
rect 79926 290898 110410 291134
rect 110646 290898 141130 291134
rect 141366 290898 171850 291134
rect 172086 290898 202570 291134
rect 202806 290898 233290 291134
rect 233526 290898 264010 291134
rect 264246 290898 294730 291134
rect 294966 290898 325450 291134
rect 325686 290898 356170 291134
rect 356406 290898 386890 291134
rect 387126 290898 417610 291134
rect 417846 290898 448330 291134
rect 448566 290898 479050 291134
rect 479286 290898 509770 291134
rect 510006 290898 540490 291134
rect 540726 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 33610 273454
rect 33846 273218 64330 273454
rect 64566 273218 95050 273454
rect 95286 273218 125770 273454
rect 126006 273218 156490 273454
rect 156726 273218 187210 273454
rect 187446 273218 217930 273454
rect 218166 273218 248650 273454
rect 248886 273218 279370 273454
rect 279606 273218 310090 273454
rect 310326 273218 340810 273454
rect 341046 273218 371530 273454
rect 371766 273218 402250 273454
rect 402486 273218 432970 273454
rect 433206 273218 463690 273454
rect 463926 273218 494410 273454
rect 494646 273218 525130 273454
rect 525366 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 33610 273134
rect 33846 272898 64330 273134
rect 64566 272898 95050 273134
rect 95286 272898 125770 273134
rect 126006 272898 156490 273134
rect 156726 272898 187210 273134
rect 187446 272898 217930 273134
rect 218166 272898 248650 273134
rect 248886 272898 279370 273134
rect 279606 272898 310090 273134
rect 310326 272898 340810 273134
rect 341046 272898 371530 273134
rect 371766 272898 402250 273134
rect 402486 272898 432970 273134
rect 433206 272898 463690 273134
rect 463926 272898 494410 273134
rect 494646 272898 525130 273134
rect 525366 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 18250 255454
rect 18486 255218 48970 255454
rect 49206 255218 79690 255454
rect 79926 255218 110410 255454
rect 110646 255218 141130 255454
rect 141366 255218 171850 255454
rect 172086 255218 202570 255454
rect 202806 255218 233290 255454
rect 233526 255218 264010 255454
rect 264246 255218 294730 255454
rect 294966 255218 325450 255454
rect 325686 255218 356170 255454
rect 356406 255218 386890 255454
rect 387126 255218 417610 255454
rect 417846 255218 448330 255454
rect 448566 255218 479050 255454
rect 479286 255218 509770 255454
rect 510006 255218 540490 255454
rect 540726 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 18250 255134
rect 18486 254898 48970 255134
rect 49206 254898 79690 255134
rect 79926 254898 110410 255134
rect 110646 254898 141130 255134
rect 141366 254898 171850 255134
rect 172086 254898 202570 255134
rect 202806 254898 233290 255134
rect 233526 254898 264010 255134
rect 264246 254898 294730 255134
rect 294966 254898 325450 255134
rect 325686 254898 356170 255134
rect 356406 254898 386890 255134
rect 387126 254898 417610 255134
rect 417846 254898 448330 255134
rect 448566 254898 479050 255134
rect 479286 254898 509770 255134
rect 510006 254898 540490 255134
rect 540726 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 33610 237454
rect 33846 237218 64330 237454
rect 64566 237218 95050 237454
rect 95286 237218 125770 237454
rect 126006 237218 156490 237454
rect 156726 237218 187210 237454
rect 187446 237218 217930 237454
rect 218166 237218 248650 237454
rect 248886 237218 279370 237454
rect 279606 237218 310090 237454
rect 310326 237218 340810 237454
rect 341046 237218 371530 237454
rect 371766 237218 402250 237454
rect 402486 237218 432970 237454
rect 433206 237218 463690 237454
rect 463926 237218 494410 237454
rect 494646 237218 525130 237454
rect 525366 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 33610 237134
rect 33846 236898 64330 237134
rect 64566 236898 95050 237134
rect 95286 236898 125770 237134
rect 126006 236898 156490 237134
rect 156726 236898 187210 237134
rect 187446 236898 217930 237134
rect 218166 236898 248650 237134
rect 248886 236898 279370 237134
rect 279606 236898 310090 237134
rect 310326 236898 340810 237134
rect 341046 236898 371530 237134
rect 371766 236898 402250 237134
rect 402486 236898 432970 237134
rect 433206 236898 463690 237134
rect 463926 236898 494410 237134
rect 494646 236898 525130 237134
rect 525366 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 18250 219454
rect 18486 219218 48970 219454
rect 49206 219218 79690 219454
rect 79926 219218 110410 219454
rect 110646 219218 141130 219454
rect 141366 219218 171850 219454
rect 172086 219218 202570 219454
rect 202806 219218 233290 219454
rect 233526 219218 264010 219454
rect 264246 219218 294730 219454
rect 294966 219218 325450 219454
rect 325686 219218 356170 219454
rect 356406 219218 386890 219454
rect 387126 219218 417610 219454
rect 417846 219218 448330 219454
rect 448566 219218 479050 219454
rect 479286 219218 509770 219454
rect 510006 219218 540490 219454
rect 540726 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 18250 219134
rect 18486 218898 48970 219134
rect 49206 218898 79690 219134
rect 79926 218898 110410 219134
rect 110646 218898 141130 219134
rect 141366 218898 171850 219134
rect 172086 218898 202570 219134
rect 202806 218898 233290 219134
rect 233526 218898 264010 219134
rect 264246 218898 294730 219134
rect 294966 218898 325450 219134
rect 325686 218898 356170 219134
rect 356406 218898 386890 219134
rect 387126 218898 417610 219134
rect 417846 218898 448330 219134
rect 448566 218898 479050 219134
rect 479286 218898 509770 219134
rect 510006 218898 540490 219134
rect 540726 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 33610 201454
rect 33846 201218 64330 201454
rect 64566 201218 95050 201454
rect 95286 201218 125770 201454
rect 126006 201218 156490 201454
rect 156726 201218 187210 201454
rect 187446 201218 217930 201454
rect 218166 201218 248650 201454
rect 248886 201218 279370 201454
rect 279606 201218 310090 201454
rect 310326 201218 340810 201454
rect 341046 201218 371530 201454
rect 371766 201218 402250 201454
rect 402486 201218 432970 201454
rect 433206 201218 463690 201454
rect 463926 201218 494410 201454
rect 494646 201218 525130 201454
rect 525366 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 33610 201134
rect 33846 200898 64330 201134
rect 64566 200898 95050 201134
rect 95286 200898 125770 201134
rect 126006 200898 156490 201134
rect 156726 200898 187210 201134
rect 187446 200898 217930 201134
rect 218166 200898 248650 201134
rect 248886 200898 279370 201134
rect 279606 200898 310090 201134
rect 310326 200898 340810 201134
rect 341046 200898 371530 201134
rect 371766 200898 402250 201134
rect 402486 200898 432970 201134
rect 433206 200898 463690 201134
rect 463926 200898 494410 201134
rect 494646 200898 525130 201134
rect 525366 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 18250 183454
rect 18486 183218 48970 183454
rect 49206 183218 79690 183454
rect 79926 183218 110410 183454
rect 110646 183218 141130 183454
rect 141366 183218 171850 183454
rect 172086 183218 202570 183454
rect 202806 183218 233290 183454
rect 233526 183218 264010 183454
rect 264246 183218 294730 183454
rect 294966 183218 325450 183454
rect 325686 183218 356170 183454
rect 356406 183218 386890 183454
rect 387126 183218 417610 183454
rect 417846 183218 448330 183454
rect 448566 183218 479050 183454
rect 479286 183218 509770 183454
rect 510006 183218 540490 183454
rect 540726 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 18250 183134
rect 18486 182898 48970 183134
rect 49206 182898 79690 183134
rect 79926 182898 110410 183134
rect 110646 182898 141130 183134
rect 141366 182898 171850 183134
rect 172086 182898 202570 183134
rect 202806 182898 233290 183134
rect 233526 182898 264010 183134
rect 264246 182898 294730 183134
rect 294966 182898 325450 183134
rect 325686 182898 356170 183134
rect 356406 182898 386890 183134
rect 387126 182898 417610 183134
rect 417846 182898 448330 183134
rect 448566 182898 479050 183134
rect 479286 182898 509770 183134
rect 510006 182898 540490 183134
rect 540726 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 33610 165454
rect 33846 165218 64330 165454
rect 64566 165218 95050 165454
rect 95286 165218 125770 165454
rect 126006 165218 156490 165454
rect 156726 165218 187210 165454
rect 187446 165218 217930 165454
rect 218166 165218 248650 165454
rect 248886 165218 279370 165454
rect 279606 165218 310090 165454
rect 310326 165218 340810 165454
rect 341046 165218 371530 165454
rect 371766 165218 402250 165454
rect 402486 165218 432970 165454
rect 433206 165218 463690 165454
rect 463926 165218 494410 165454
rect 494646 165218 525130 165454
rect 525366 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 33610 165134
rect 33846 164898 64330 165134
rect 64566 164898 95050 165134
rect 95286 164898 125770 165134
rect 126006 164898 156490 165134
rect 156726 164898 187210 165134
rect 187446 164898 217930 165134
rect 218166 164898 248650 165134
rect 248886 164898 279370 165134
rect 279606 164898 310090 165134
rect 310326 164898 340810 165134
rect 341046 164898 371530 165134
rect 371766 164898 402250 165134
rect 402486 164898 432970 165134
rect 433206 164898 463690 165134
rect 463926 164898 494410 165134
rect 494646 164898 525130 165134
rect 525366 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 18250 147454
rect 18486 147218 48970 147454
rect 49206 147218 79690 147454
rect 79926 147218 110410 147454
rect 110646 147218 141130 147454
rect 141366 147218 171850 147454
rect 172086 147218 202570 147454
rect 202806 147218 233290 147454
rect 233526 147218 264010 147454
rect 264246 147218 294730 147454
rect 294966 147218 325450 147454
rect 325686 147218 356170 147454
rect 356406 147218 386890 147454
rect 387126 147218 417610 147454
rect 417846 147218 448330 147454
rect 448566 147218 479050 147454
rect 479286 147218 509770 147454
rect 510006 147218 540490 147454
rect 540726 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 18250 147134
rect 18486 146898 48970 147134
rect 49206 146898 79690 147134
rect 79926 146898 110410 147134
rect 110646 146898 141130 147134
rect 141366 146898 171850 147134
rect 172086 146898 202570 147134
rect 202806 146898 233290 147134
rect 233526 146898 264010 147134
rect 264246 146898 294730 147134
rect 294966 146898 325450 147134
rect 325686 146898 356170 147134
rect 356406 146898 386890 147134
rect 387126 146898 417610 147134
rect 417846 146898 448330 147134
rect 448566 146898 479050 147134
rect 479286 146898 509770 147134
rect 510006 146898 540490 147134
rect 540726 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 33610 129454
rect 33846 129218 64330 129454
rect 64566 129218 95050 129454
rect 95286 129218 125770 129454
rect 126006 129218 156490 129454
rect 156726 129218 187210 129454
rect 187446 129218 217930 129454
rect 218166 129218 248650 129454
rect 248886 129218 279370 129454
rect 279606 129218 310090 129454
rect 310326 129218 340810 129454
rect 341046 129218 371530 129454
rect 371766 129218 402250 129454
rect 402486 129218 432970 129454
rect 433206 129218 463690 129454
rect 463926 129218 494410 129454
rect 494646 129218 525130 129454
rect 525366 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 33610 129134
rect 33846 128898 64330 129134
rect 64566 128898 95050 129134
rect 95286 128898 125770 129134
rect 126006 128898 156490 129134
rect 156726 128898 187210 129134
rect 187446 128898 217930 129134
rect 218166 128898 248650 129134
rect 248886 128898 279370 129134
rect 279606 128898 310090 129134
rect 310326 128898 340810 129134
rect 341046 128898 371530 129134
rect 371766 128898 402250 129134
rect 402486 128898 432970 129134
rect 433206 128898 463690 129134
rect 463926 128898 494410 129134
rect 494646 128898 525130 129134
rect 525366 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 18250 111454
rect 18486 111218 48970 111454
rect 49206 111218 79690 111454
rect 79926 111218 110410 111454
rect 110646 111218 141130 111454
rect 141366 111218 171850 111454
rect 172086 111218 202570 111454
rect 202806 111218 233290 111454
rect 233526 111218 264010 111454
rect 264246 111218 294730 111454
rect 294966 111218 325450 111454
rect 325686 111218 356170 111454
rect 356406 111218 386890 111454
rect 387126 111218 417610 111454
rect 417846 111218 448330 111454
rect 448566 111218 479050 111454
rect 479286 111218 509770 111454
rect 510006 111218 540490 111454
rect 540726 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 18250 111134
rect 18486 110898 48970 111134
rect 49206 110898 79690 111134
rect 79926 110898 110410 111134
rect 110646 110898 141130 111134
rect 141366 110898 171850 111134
rect 172086 110898 202570 111134
rect 202806 110898 233290 111134
rect 233526 110898 264010 111134
rect 264246 110898 294730 111134
rect 294966 110898 325450 111134
rect 325686 110898 356170 111134
rect 356406 110898 386890 111134
rect 387126 110898 417610 111134
rect 417846 110898 448330 111134
rect 448566 110898 479050 111134
rect 479286 110898 509770 111134
rect 510006 110898 540490 111134
rect 540726 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 33610 93454
rect 33846 93218 64330 93454
rect 64566 93218 95050 93454
rect 95286 93218 125770 93454
rect 126006 93218 156490 93454
rect 156726 93218 187210 93454
rect 187446 93218 217930 93454
rect 218166 93218 248650 93454
rect 248886 93218 279370 93454
rect 279606 93218 310090 93454
rect 310326 93218 340810 93454
rect 341046 93218 371530 93454
rect 371766 93218 402250 93454
rect 402486 93218 432970 93454
rect 433206 93218 463690 93454
rect 463926 93218 494410 93454
rect 494646 93218 525130 93454
rect 525366 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 33610 93134
rect 33846 92898 64330 93134
rect 64566 92898 95050 93134
rect 95286 92898 125770 93134
rect 126006 92898 156490 93134
rect 156726 92898 187210 93134
rect 187446 92898 217930 93134
rect 218166 92898 248650 93134
rect 248886 92898 279370 93134
rect 279606 92898 310090 93134
rect 310326 92898 340810 93134
rect 341046 92898 371530 93134
rect 371766 92898 402250 93134
rect 402486 92898 432970 93134
rect 433206 92898 463690 93134
rect 463926 92898 494410 93134
rect 494646 92898 525130 93134
rect 525366 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 18250 75454
rect 18486 75218 48970 75454
rect 49206 75218 79690 75454
rect 79926 75218 110410 75454
rect 110646 75218 141130 75454
rect 141366 75218 171850 75454
rect 172086 75218 202570 75454
rect 202806 75218 233290 75454
rect 233526 75218 264010 75454
rect 264246 75218 294730 75454
rect 294966 75218 325450 75454
rect 325686 75218 356170 75454
rect 356406 75218 386890 75454
rect 387126 75218 417610 75454
rect 417846 75218 448330 75454
rect 448566 75218 479050 75454
rect 479286 75218 509770 75454
rect 510006 75218 540490 75454
rect 540726 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 18250 75134
rect 18486 74898 48970 75134
rect 49206 74898 79690 75134
rect 79926 74898 110410 75134
rect 110646 74898 141130 75134
rect 141366 74898 171850 75134
rect 172086 74898 202570 75134
rect 202806 74898 233290 75134
rect 233526 74898 264010 75134
rect 264246 74898 294730 75134
rect 294966 74898 325450 75134
rect 325686 74898 356170 75134
rect 356406 74898 386890 75134
rect 387126 74898 417610 75134
rect 417846 74898 448330 75134
rect 448566 74898 479050 75134
rect 479286 74898 509770 75134
rect 510006 74898 540490 75134
rect 540726 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 33610 57454
rect 33846 57218 64330 57454
rect 64566 57218 95050 57454
rect 95286 57218 125770 57454
rect 126006 57218 156490 57454
rect 156726 57218 187210 57454
rect 187446 57218 217930 57454
rect 218166 57218 248650 57454
rect 248886 57218 279370 57454
rect 279606 57218 310090 57454
rect 310326 57218 340810 57454
rect 341046 57218 371530 57454
rect 371766 57218 402250 57454
rect 402486 57218 432970 57454
rect 433206 57218 463690 57454
rect 463926 57218 494410 57454
rect 494646 57218 525130 57454
rect 525366 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 33610 57134
rect 33846 56898 64330 57134
rect 64566 56898 95050 57134
rect 95286 56898 125770 57134
rect 126006 56898 156490 57134
rect 156726 56898 187210 57134
rect 187446 56898 217930 57134
rect 218166 56898 248650 57134
rect 248886 56898 279370 57134
rect 279606 56898 310090 57134
rect 310326 56898 340810 57134
rect 341046 56898 371530 57134
rect 371766 56898 402250 57134
rect 402486 56898 432970 57134
rect 433206 56898 463690 57134
rect 463926 56898 494410 57134
rect 494646 56898 525130 57134
rect 525366 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 1640738188
transform 1 0 14000 0 1 50000
box 0 0 539474 620000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 672000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 672000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 672000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 672000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 672000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 672000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 672000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 672000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 672000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 672000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 672000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 672000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 672000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 672000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 672000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 672000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 672000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 672000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 672000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 672000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 672000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 672000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 672000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 672000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 672000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 672000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 672000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 672000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 672000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 672000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 672000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 672000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 672000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 672000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 672000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 672000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 672000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 672000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 672000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 672000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 672000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 672000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 672000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 672000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 672000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 672000 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 672000 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 672000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 672000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 672000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 672000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 672000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 672000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 672000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 672000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 672000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 672000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 672000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 672000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 672000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 672000 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 672000 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 672000 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 672000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 672000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 672000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 672000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 672000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 672000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 672000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 672000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 672000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 672000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 672000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 672000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 672000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 672000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 672000 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 672000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 672000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 672000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 672000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 672000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 672000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 672000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 672000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 672000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 672000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 672000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 672000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 672000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 672000 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 672000 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 672000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 672000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 672000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 672000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 672000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 672000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 672000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 672000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 672000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 672000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 672000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 672000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 672000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 672000 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 672000 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 672000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 672000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 672000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 672000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 672000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 672000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 672000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 672000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 672000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 672000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 672000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 672000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 672000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
